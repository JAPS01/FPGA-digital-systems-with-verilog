`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:31:35 04/29/2021 
// Design Name: 
// Module Name:    Personaje 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Personaje(
input enable,
input clock,
input [9:0] X, Y,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg imagen);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= X & hcount < X + RESOLUCION_X & vcount >= Y & vcount < Y + RESOLUCION_Y)
		begin
			if (Batman[vcount - Y][hcount - X][8] == 1'b1)
			begin
				red   <= Batman[vcount- Y][hcount- X][7:5];
				green <= Batman[vcount- Y][hcount- X][4:2];
            blue 	<= Batman[vcount- Y][hcount- X][1:0];
				imagen  <= 1'b1;
			end
			else
				imagen <= 0;
			end
		else
		imagen <= 0;
	end
end

parameter RESOLUCION_X = 40;
parameter RESOLUCION_Y = 40;
wire [8:0] Batman[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign Batman[1][18] = 9'b100000000;
assign Batman[1][25] = 9'b100000000;
assign Batman[1][26] = 9'b100000000;
assign Batman[2][17] = 9'b100000000;
assign Batman[2][18] = 9'b100000000;
assign Batman[2][19] = 9'b100000000;
assign Batman[2][21] = 9'b100000000;
assign Batman[2][22] = 9'b100000000;
assign Batman[2][23] = 9'b100000000;
assign Batman[2][25] = 9'b100000000;
assign Batman[2][26] = 9'b100000000;
assign Batman[3][17] = 9'b100000000;
assign Batman[3][18] = 9'b100100100;
assign Batman[3][19] = 9'b100000000;
assign Batman[3][20] = 9'b100000000;
assign Batman[3][21] = 9'b100100100;
assign Batman[3][22] = 9'b100100100;
assign Batman[3][23] = 9'b100100100;
assign Batman[3][24] = 9'b100000000;
assign Batman[3][25] = 9'b100000000;
assign Batman[3][26] = 9'b100000000;
assign Batman[4][17] = 9'b100000000;
assign Batman[4][18] = 9'b100100100;
assign Batman[4][19] = 9'b100000000;
assign Batman[4][20] = 9'b100100100;
assign Batman[4][21] = 9'b100100100;
assign Batman[4][22] = 9'b101001001;
assign Batman[4][23] = 9'b101101101;
assign Batman[4][24] = 9'b101001001;
assign Batman[4][25] = 9'b100100100;
assign Batman[4][26] = 9'b100000000;
assign Batman[5][17] = 9'b100000000;
assign Batman[5][18] = 9'b100100100;
assign Batman[5][19] = 9'b100100100;
assign Batman[5][20] = 9'b100100100;
assign Batman[5][21] = 9'b101001001;
assign Batman[5][22] = 9'b101101101;
assign Batman[5][23] = 9'b101101101;
assign Batman[5][24] = 9'b101101101;
assign Batman[5][25] = 9'b101001001;
assign Batman[5][26] = 9'b100000000;
assign Batman[6][16] = 9'b100000000;
assign Batman[6][17] = 9'b100000000;
assign Batman[6][18] = 9'b100100100;
assign Batman[6][19] = 9'b100100100;
assign Batman[6][20] = 9'b100100100;
assign Batman[6][21] = 9'b101101101;
assign Batman[6][22] = 9'b101101101;
assign Batman[6][23] = 9'b101101101;
assign Batman[6][24] = 9'b101101101;
assign Batman[6][25] = 9'b101101101;
assign Batman[6][26] = 9'b100100100;
assign Batman[6][27] = 9'b100000000;
assign Batman[7][16] = 9'b100000000;
assign Batman[7][17] = 9'b100000000;
assign Batman[7][18] = 9'b100000000;
assign Batman[7][19] = 9'b100100100;
assign Batman[7][20] = 9'b100100100;
assign Batman[7][21] = 9'b101001001;
assign Batman[7][22] = 9'b101101101;
assign Batman[7][23] = 9'b101101101;
assign Batman[7][24] = 9'b101101101;
assign Batman[7][25] = 9'b101101101;
assign Batman[7][26] = 9'b101101101;
assign Batman[7][27] = 9'b100000000;
assign Batman[8][16] = 9'b100000000;
assign Batman[8][17] = 9'b100000000;
assign Batman[8][18] = 9'b100000000;
assign Batman[8][19] = 9'b100000000;
assign Batman[8][20] = 9'b100000000;
assign Batman[8][21] = 9'b100000000;
assign Batman[8][22] = 9'b101001001;
assign Batman[8][23] = 9'b101101101;
assign Batman[8][24] = 9'b101101101;
assign Batman[8][25] = 9'b101101101;
assign Batman[8][26] = 9'b101101101;
assign Batman[8][27] = 9'b100000000;
assign Batman[9][16] = 9'b100000000;
assign Batman[9][17] = 9'b100000000;
assign Batman[9][18] = 9'b100000000;
assign Batman[9][19] = 9'b100000000;
assign Batman[9][20] = 9'b100000000;
assign Batman[9][22] = 9'b100000000;
assign Batman[9][23] = 9'b100100100;
assign Batman[9][24] = 9'b101101101;
assign Batman[9][25] = 9'b101101101;
assign Batman[9][26] = 9'b101001001;
assign Batman[9][27] = 9'b100000000;
assign Batman[10][17] = 9'b100000000;
assign Batman[10][18] = 9'b100000000;
assign Batman[10][19] = 9'b100000000;
assign Batman[10][20] = 9'b100000000;
assign Batman[10][21] = 9'b100000000;
assign Batman[10][23] = 9'b100000000;
assign Batman[10][24] = 9'b100100100;
assign Batman[10][25] = 9'b101001001;
assign Batman[10][26] = 9'b100100100;
assign Batman[10][27] = 9'b100000000;
assign Batman[11][17] = 9'b100000000;
assign Batman[11][18] = 9'b100000000;
assign Batman[11][19] = 9'b100000000;
assign Batman[11][20] = 9'b100100100;
assign Batman[11][21] = 9'b100000000;
assign Batman[11][22] = 9'b100000000;
assign Batman[11][23] = 9'b100000000;
assign Batman[11][24] = 9'b100000000;
assign Batman[11][25] = 9'b101001000;
assign Batman[11][26] = 9'b100100100;
assign Batman[12][17] = 9'b100000000;
assign Batman[12][18] = 9'b100000000;
assign Batman[12][19] = 9'b100000000;
assign Batman[12][20] = 9'b100100100;
assign Batman[12][21] = 9'b110001101;
assign Batman[12][22] = 9'b110001101;
assign Batman[12][23] = 9'b101101000;
assign Batman[12][24] = 9'b110001101;
assign Batman[12][25] = 9'b110101101;
assign Batman[12][26] = 9'b100100100;
assign Batman[13][17] = 9'b100000000;
assign Batman[13][18] = 9'b100100100;
assign Batman[13][19] = 9'b100100100;
assign Batman[13][20] = 9'b100100100;
assign Batman[13][21] = 9'b110101101;
assign Batman[13][22] = 9'b110001101;
assign Batman[13][23] = 9'b101001000;
assign Batman[13][24] = 9'b100100100;
assign Batman[13][25] = 9'b100100100;
assign Batman[14][15] = 9'b100000000;
assign Batman[14][16] = 9'b100000000;
assign Batman[14][17] = 9'b100100100;
assign Batman[14][18] = 9'b100100100;
assign Batman[14][19] = 9'b101001000;
assign Batman[14][20] = 9'b100000000;
assign Batman[14][21] = 9'b100100100;
assign Batman[14][22] = 9'b101001000;
assign Batman[14][23] = 9'b101001000;
assign Batman[14][24] = 9'b100100100;
assign Batman[15][14] = 9'b100000000;
assign Batman[15][15] = 9'b100100100;
assign Batman[15][16] = 9'b101001000;
assign Batman[15][17] = 9'b101001001;
assign Batman[15][19] = 9'b100000000;
assign Batman[15][20] = 9'b100000000;
assign Batman[15][21] = 9'b100000000;
assign Batman[15][22] = 9'b100000000;
assign Batman[15][23] = 9'b100000000;
assign Batman[15][24] = 9'b100000000;
assign Batman[15][25] = 9'b100000000;
assign Batman[15][26] = 9'b100000000;
assign Batman[16][13] = 9'b100000000;
assign Batman[16][14] = 9'b100100100;
assign Batman[16][15] = 9'b110010010;
assign Batman[16][17] = 9'b100000000;
assign Batman[16][18] = 9'b101001001;
assign Batman[16][19] = 9'b101001000;
assign Batman[16][21] = 9'b100000000;
assign Batman[16][22] = 9'b100000000;
assign Batman[16][23] = 9'b100000000;
assign Batman[16][24] = 9'b100000000;
assign Batman[16][25] = 9'b100000000;
assign Batman[16][26] = 9'b100000000;
assign Batman[17][13] = 9'b100000000;
assign Batman[17][14] = 9'b101001000;
assign Batman[17][15] = 9'b101001001;
assign Batman[17][16] = 9'b101101101;
assign Batman[17][17] = 9'b100100100;
assign Batman[17][18] = 9'b100100100;
assign Batman[17][19] = 9'b101001001;
assign Batman[17][20] = 9'b101001000;
assign Batman[17][21] = 9'b100000000;
assign Batman[17][22] = 9'b100000000;
assign Batman[17][23] = 9'b100100100;
assign Batman[17][24] = 9'b100000000;
assign Batman[17][25] = 9'b100000000;
assign Batman[17][26] = 9'b100000000;
assign Batman[18][13] = 9'b100000000;
assign Batman[18][14] = 9'b101001001;
assign Batman[18][15] = 9'b101001000;
assign Batman[18][16] = 9'b100100100;
assign Batman[18][17] = 9'b101001000;
assign Batman[18][19] = 9'b100100100;
assign Batman[18][20] = 9'b101101101;
assign Batman[18][21] = 9'b101101101;
assign Batman[18][22] = 9'b101001000;
assign Batman[18][23] = 9'b100000000;
assign Batman[18][24] = 9'b100100100;
assign Batman[18][25] = 9'b100100100;
assign Batman[18][26] = 9'b100000000;
assign Batman[18][27] = 9'b100000000;
assign Batman[19][12] = 9'b100000000;
assign Batman[19][13] = 9'b100000000;
assign Batman[19][14] = 9'b100100100;
assign Batman[19][15] = 9'b101001001;
assign Batman[19][16] = 9'b100100100;
assign Batman[19][17] = 9'b100000000;
assign Batman[19][18] = 9'b100100100;
assign Batman[19][19] = 9'b101101101;
assign Batman[19][20] = 9'b100100100;
assign Batman[19][21] = 9'b101001000;
assign Batman[19][22] = 9'b101001000;
assign Batman[19][23] = 9'b100100100;
assign Batman[19][24] = 9'b101001001;
assign Batman[19][25] = 9'b100100100;
assign Batman[19][26] = 9'b100000000;
assign Batman[19][27] = 9'b100000000;
assign Batman[20][12] = 9'b100000000;
assign Batman[20][13] = 9'b101001001;
assign Batman[20][14] = 9'b101001001;
assign Batman[20][16] = 9'b100000000;
assign Batman[20][17] = 9'b100000000;
assign Batman[20][18] = 9'b100000000;
assign Batman[20][19] = 9'b100100100;
assign Batman[20][21] = 9'b100100100;
assign Batman[20][22] = 9'b101101101;
assign Batman[20][23] = 9'b101001000;
assign Batman[20][25] = 9'b100000000;
assign Batman[20][26] = 9'b100000000;
assign Batman[20][27] = 9'b100000000;
assign Batman[21][11] = 9'b100000000;
assign Batman[21][12] = 9'b100000000;
assign Batman[21][13] = 9'b100100100;
assign Batman[21][14] = 9'b100100100;
assign Batman[21][15] = 9'b100000000;
assign Batman[21][16] = 9'b100000000;
assign Batman[21][17] = 9'b100100100;
assign Batman[21][18] = 9'b100100100;
assign Batman[21][19] = 9'b100000000;
assign Batman[21][20] = 9'b100000000;
assign Batman[21][21] = 9'b100000000;
assign Batman[21][22] = 9'b100000000;
assign Batman[21][23] = 9'b100000000;
assign Batman[21][24] = 9'b100000000;
assign Batman[21][25] = 9'b100000000;
assign Batman[21][26] = 9'b100000000;
assign Batman[21][27] = 9'b100000000;
assign Batman[22][11] = 9'b100000000;
assign Batman[22][12] = 9'b100000000;
assign Batman[22][13] = 9'b100000000;
assign Batman[22][14] = 9'b100000000;
assign Batman[22][15] = 9'b100000000;
assign Batman[22][16] = 9'b100000000;
assign Batman[22][17] = 9'b100100100;
assign Batman[22][18] = 9'b100100100;
assign Batman[22][19] = 9'b100000000;
assign Batman[22][20] = 9'b101000100;
assign Batman[22][21] = 9'b101000100;
assign Batman[22][22] = 9'b101000100;
assign Batman[22][23] = 9'b101000100;
assign Batman[22][24] = 9'b101101000;
assign Batman[22][25] = 9'b100100100;
assign Batman[22][26] = 9'b100000000;
assign Batman[22][27] = 9'b100000000;
assign Batman[23][10] = 9'b100000000;
assign Batman[23][11] = 9'b100000000;
assign Batman[23][12] = 9'b100000000;
assign Batman[23][13] = 9'b100100100;
assign Batman[23][14] = 9'b100100100;
assign Batman[23][15] = 9'b100000000;
assign Batman[23][16] = 9'b100000000;
assign Batman[23][17] = 9'b100100100;
assign Batman[23][18] = 9'b100000000;
assign Batman[23][19] = 9'b101000100;
assign Batman[23][20] = 9'b110101100;
assign Batman[23][21] = 9'b111110000;
assign Batman[23][22] = 9'b110101100;
assign Batman[23][23] = 9'b110101100;
assign Batman[23][24] = 9'b111110001;
assign Batman[23][25] = 9'b101000100;
assign Batman[23][26] = 9'b100000000;
assign Batman[23][27] = 9'b100000000;
assign Batman[24][10] = 9'b100000000;
assign Batman[24][11] = 9'b100100100;
assign Batman[24][12] = 9'b100000000;
assign Batman[24][13] = 9'b100100100;
assign Batman[24][14] = 9'b101001000;
assign Batman[24][15] = 9'b100100100;
assign Batman[24][16] = 9'b100000000;
assign Batman[24][17] = 9'b100000000;
assign Batman[24][18] = 9'b100000000;
assign Batman[24][19] = 9'b100000000;
assign Batman[24][20] = 9'b100000000;
assign Batman[24][21] = 9'b100000000;
assign Batman[24][22] = 9'b100000000;
assign Batman[24][23] = 9'b100000000;
assign Batman[24][24] = 9'b100000000;
assign Batman[24][25] = 9'b100000000;
assign Batman[24][26] = 9'b100000000;
assign Batman[24][27] = 9'b100000000;
assign Batman[24][28] = 9'b100000000;
assign Batman[25][9] = 9'b100000000;
assign Batman[25][10] = 9'b100000000;
assign Batman[25][11] = 9'b100100100;
assign Batman[25][12] = 9'b100000000;
assign Batman[25][13] = 9'b100100100;
assign Batman[25][15] = 9'b100100100;
assign Batman[25][16] = 9'b100100100;
assign Batman[25][17] = 9'b100000000;
assign Batman[25][18] = 9'b101001001;
assign Batman[25][19] = 9'b110010010;
assign Batman[25][20] = 9'b100000000;
assign Batman[25][21] = 9'b100000000;
assign Batman[25][22] = 9'b101001000;
assign Batman[25][23] = 9'b100100100;
assign Batman[25][24] = 9'b100000000;
assign Batman[25][25] = 9'b100000000;
assign Batman[25][26] = 9'b100000000;
assign Batman[25][27] = 9'b100000000;
assign Batman[25][28] = 9'b100000000;
assign Batman[26][9] = 9'b100000000;
assign Batman[26][10] = 9'b100100100;
assign Batman[26][11] = 9'b100000000;
assign Batman[26][12] = 9'b100000000;
assign Batman[26][13] = 9'b100000000;
assign Batman[26][14] = 9'b100100100;
assign Batman[26][15] = 9'b100000000;
assign Batman[26][16] = 9'b100000000;
assign Batman[26][17] = 9'b100000000;
assign Batman[26][18] = 9'b111111111;
assign Batman[26][19] = 9'b110110110;
assign Batman[26][21] = 9'b100000000;
assign Batman[26][22] = 9'b100000000;
assign Batman[26][23] = 9'b100000000;
assign Batman[26][24] = 9'b100000000;
assign Batman[26][26] = 9'b100000000;
assign Batman[26][27] = 9'b100000000;
assign Batman[26][28] = 9'b100000000;
assign Batman[27][9] = 9'b100000000;
assign Batman[27][10] = 9'b100000000;
assign Batman[27][11] = 9'b100000000;
assign Batman[27][12] = 9'b100000000;
assign Batman[27][13] = 9'b100000000;
assign Batman[27][14] = 9'b100000000;
assign Batman[27][15] = 9'b100000000;
assign Batman[27][16] = 9'b100000000;
assign Batman[27][17] = 9'b100000000;
assign Batman[27][18] = 9'b101001001;
assign Batman[27][19] = 9'b110010010;
assign Batman[27][20] = 9'b101101101;
assign Batman[27][21] = 9'b100100100;
assign Batman[27][22] = 9'b100000000;
assign Batman[27][23] = 9'b100000000;
assign Batman[27][24] = 9'b111111111;
assign Batman[27][26] = 9'b100000000;
assign Batman[27][27] = 9'b100000000;
assign Batman[27][28] = 9'b100000000;
assign Batman[27][29] = 9'b100000000;
assign Batman[28][9] = 9'b100000000;
assign Batman[28][10] = 9'b100000000;
assign Batman[28][11] = 9'b100000000;
assign Batman[28][12] = 9'b100100100;
assign Batman[28][13] = 9'b100100100;
assign Batman[28][14] = 9'b100000000;
assign Batman[28][15] = 9'b100000000;
assign Batman[28][16] = 9'b100000000;
assign Batman[28][17] = 9'b101001000;
assign Batman[28][18] = 9'b101001001;
assign Batman[28][19] = 9'b101101101;
assign Batman[28][20] = 9'b100100100;
assign Batman[28][21] = 9'b100000000;
assign Batman[28][22] = 9'b100000000;
assign Batman[28][24] = 9'b101001000;
assign Batman[28][26] = 9'b100000000;
assign Batman[28][27] = 9'b100000000;
assign Batman[28][28] = 9'b100100100;
assign Batman[28][29] = 9'b100000000;
assign Batman[28][30] = 9'b100000000;
assign Batman[29][8] = 9'b100000000;
assign Batman[29][9] = 9'b100100100;
assign Batman[29][10] = 9'b100000000;
assign Batman[29][11] = 9'b100000000;
assign Batman[29][12] = 9'b100100100;
assign Batman[29][13] = 9'b101001001;
assign Batman[29][14] = 9'b101101101;
assign Batman[29][15] = 9'b101001001;
assign Batman[29][16] = 9'b100000000;
assign Batman[29][17] = 9'b101101101;
assign Batman[29][18] = 9'b101001001;
assign Batman[29][19] = 9'b101001000;
assign Batman[29][20] = 9'b100100100;
assign Batman[29][21] = 9'b100000000;
assign Batman[29][22] = 9'b100000000;
assign Batman[29][23] = 9'b100100100;
assign Batman[29][24] = 9'b101101101;
assign Batman[29][25] = 9'b100100100;
assign Batman[29][26] = 9'b100000000;
assign Batman[29][27] = 9'b100000000;
assign Batman[29][28] = 9'b100100100;
assign Batman[29][29] = 9'b100000000;
assign Batman[29][30] = 9'b100000000;
assign Batman[30][8] = 9'b100000000;
assign Batman[30][9] = 9'b100000000;
assign Batman[30][10] = 9'b100000000;
assign Batman[30][11] = 9'b100100100;
assign Batman[30][12] = 9'b100100100;
assign Batman[30][13] = 9'b101101101;
assign Batman[30][14] = 9'b101101101;
assign Batman[30][15] = 9'b100100100;
assign Batman[30][16] = 9'b100100100;
assign Batman[30][17] = 9'b110010001;
assign Batman[30][19] = 9'b101101101;
assign Batman[30][20] = 9'b100100100;
assign Batman[30][21] = 9'b100000000;
assign Batman[30][22] = 9'b100000000;
assign Batman[30][23] = 9'b100100100;
assign Batman[30][24] = 9'b101101101;
assign Batman[30][26] = 9'b100000000;
assign Batman[30][27] = 9'b100000000;
assign Batman[30][28] = 9'b100100100;
assign Batman[30][29] = 9'b100100100;
assign Batman[30][30] = 9'b100000000;
assign Batman[31][8] = 9'b100000000;
assign Batman[31][9] = 9'b100000000;
assign Batman[31][10] = 9'b100000000;
assign Batman[31][11] = 9'b100100100;
assign Batman[31][12] = 9'b100100100;
assign Batman[31][13] = 9'b101001001;
assign Batman[31][14] = 9'b101001001;
assign Batman[31][15] = 9'b100000000;
assign Batman[31][16] = 9'b101101101;
assign Batman[31][17] = 9'b111111111;
assign Batman[31][19] = 9'b101001001;
assign Batman[31][20] = 9'b100000000;
assign Batman[31][21] = 9'b100100100;
assign Batman[31][22] = 9'b100000000;
assign Batman[31][23] = 9'b100000000;
assign Batman[31][26] = 9'b100000000;
assign Batman[31][27] = 9'b100000000;
assign Batman[31][28] = 9'b100100100;
assign Batman[31][29] = 9'b101001001;
assign Batman[31][30] = 9'b100000000;
assign Batman[31][31] = 9'b100000000;
assign Batman[32][8] = 9'b100000000;
assign Batman[32][9] = 9'b100000000;
assign Batman[32][10] = 9'b100000000;
assign Batman[32][11] = 9'b100000000;
assign Batman[32][12] = 9'b100100100;
assign Batman[32][13] = 9'b100100100;
assign Batman[32][14] = 9'b100100100;
assign Batman[32][15] = 9'b100000000;
assign Batman[32][16] = 9'b101001001;
assign Batman[32][19] = 9'b100000000;
assign Batman[32][20] = 9'b100000000;
assign Batman[32][21] = 9'b100100100;
assign Batman[32][22] = 9'b100000000;
assign Batman[32][23] = 9'b100000000;
assign Batman[32][24] = 9'b101001000;
assign Batman[32][26] = 9'b100000000;
assign Batman[32][27] = 9'b100000000;
assign Batman[32][28] = 9'b100000000;
assign Batman[32][29] = 9'b101001000;
assign Batman[32][30] = 9'b100000000;
assign Batman[33][8] = 9'b100000000;
assign Batman[33][9] = 9'b100100100;
assign Batman[33][10] = 9'b100000000;
assign Batman[33][11] = 9'b100000000;
assign Batman[33][12] = 9'b100000000;
assign Batman[33][13] = 9'b100000000;
assign Batman[33][14] = 9'b100000000;
assign Batman[33][15] = 9'b100000000;
assign Batman[33][16] = 9'b100000000;
assign Batman[33][17] = 9'b100000100;
assign Batman[33][18] = 9'b100100100;
assign Batman[33][19] = 9'b100000000;
assign Batman[33][20] = 9'b100000000;
assign Batman[33][21] = 9'b100100100;
assign Batman[33][22] = 9'b100000000;
assign Batman[33][23] = 9'b100000000;
assign Batman[33][24] = 9'b100000000;
assign Batman[33][25] = 9'b100100100;
assign Batman[33][26] = 9'b100000000;
assign Batman[33][27] = 9'b100000000;
assign Batman[33][28] = 9'b100000000;
assign Batman[33][29] = 9'b100000000;
assign Batman[33][30] = 9'b100000000;
assign Batman[34][8] = 9'b100000000;
assign Batman[34][9] = 9'b100100100;
assign Batman[34][10] = 9'b100000000;
assign Batman[34][12] = 9'b100000000;
assign Batman[34][13] = 9'b100000000;
assign Batman[34][14] = 9'b100000000;
assign Batman[34][15] = 9'b100000000;
assign Batman[34][16] = 9'b100100100;
assign Batman[34][17] = 9'b100100100;
assign Batman[34][18] = 9'b100000000;
assign Batman[34][19] = 9'b100000000;
assign Batman[34][20] = 9'b100000000;
assign Batman[34][21] = 9'b100000000;
assign Batman[34][22] = 9'b100000000;
assign Batman[34][23] = 9'b100000000;
assign Batman[34][24] = 9'b100100100;
assign Batman[34][25] = 9'b100100100;
assign Batman[34][26] = 9'b100000000;
assign Batman[34][29] = 9'b100000000;
assign Batman[34][30] = 9'b100000000;
assign Batman[35][8] = 9'b100000000;
assign Batman[35][9] = 9'b100000000;
assign Batman[35][10] = 9'b100000000;
assign Batman[35][13] = 9'b100000000;
assign Batman[35][14] = 9'b100000000;
assign Batman[35][15] = 9'b100100100;
assign Batman[35][16] = 9'b101101101;
assign Batman[35][17] = 9'b101001001;
assign Batman[35][18] = 9'b100000000;
assign Batman[35][22] = 9'b100000000;
assign Batman[35][23] = 9'b100000000;
assign Batman[35][24] = 9'b100100100;
assign Batman[35][26] = 9'b100100100;
assign Batman[35][27] = 9'b100000000;
assign Batman[36][13] = 9'b100000000;
assign Batman[36][14] = 9'b100000000;
assign Batman[36][15] = 9'b100100100;
assign Batman[36][16] = 9'b101001001;
assign Batman[36][17] = 9'b100000000;
assign Batman[36][18] = 9'b100000000;
assign Batman[36][23] = 9'b100000000;
assign Batman[36][24] = 9'b100000000;
assign Batman[36][25] = 9'b100100100;
assign Batman[36][26] = 9'b100100100;
assign Batman[36][27] = 9'b100000000;
assign Batman[36][28] = 9'b100000000;
assign Batman[37][13] = 9'b100000000;
assign Batman[37][14] = 9'b100000000;
assign Batman[37][15] = 9'b100000000;
assign Batman[37][16] = 9'b100000000;
assign Batman[37][17] = 9'b100000000;
assign Batman[37][18] = 9'b100000000;
assign Batman[37][24] = 9'b100000000;
assign Batman[37][25] = 9'b100000000;
assign Batman[37][26] = 9'b100000000;
assign Batman[37][27] = 9'b100000000;
assign Batman[37][28] = 9'b100000000;
assign Batman[38][14] = 9'b100000000;
assign Batman[38][15] = 9'b100000000;
assign Batman[38][16] = 9'b100000000;
assign Batman[38][17] = 9'b100000000;
//Total de Lineas = 535


endmodule

