`timescale 1ns / 1ps

module Logo(
input enable,
input clock,
input [9:0] X, Y,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg imagen);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= X & hcount < X + RESOLUCION_X & vcount >= Y & vcount < Y + RESOLUCION_Y)
		begin
			if (Simbolo[vcount - Y][hcount - X][8] == 1'b1)
			begin
				red   <= Simbolo[vcount- Y][hcount- X][7:5];
				green <= Simbolo[vcount- Y][hcount- X][4:2];
            blue 	<= Simbolo[vcount- Y][hcount- X][1:0];
				imagen  <= 1'b1;
			end
			else
				imagen <= 0;
			end
		else
		imagen <= 0;
	end
end

parameter RESOLUCION_X = 70;
parameter RESOLUCION_Y = 40;
wire [8:0] Simbolo[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign Simbolo[9][20] = 9'b100100000;
assign Simbolo[9][21] = 9'b100100000;
assign Simbolo[9][22] = 9'b101100100;
assign Simbolo[9][23] = 9'b111110001;
assign Simbolo[9][31] = 9'b100000000;
assign Simbolo[9][32] = 9'b100000000;
assign Simbolo[9][37] = 9'b100000000;
assign Simbolo[9][38] = 9'b100000000;
assign Simbolo[9][47] = 9'b101100100;
assign Simbolo[9][48] = 9'b100100000;
assign Simbolo[9][49] = 9'b100100000;
assign Simbolo[10][17] = 9'b100000000;
assign Simbolo[10][18] = 9'b100000000;
assign Simbolo[10][19] = 9'b100000000;
assign Simbolo[10][20] = 9'b100000000;
assign Simbolo[10][21] = 9'b101000100;
assign Simbolo[10][22] = 9'b111110001;
assign Simbolo[10][31] = 9'b100000000;
assign Simbolo[10][32] = 9'b100000000;
assign Simbolo[10][33] = 9'b100000000;
assign Simbolo[10][34] = 9'b100000000;
assign Simbolo[10][35] = 9'b100000000;
assign Simbolo[10][36] = 9'b100000000;
assign Simbolo[10][37] = 9'b100000000;
assign Simbolo[10][38] = 9'b100000000;
assign Simbolo[10][47] = 9'b111110001;
assign Simbolo[10][48] = 9'b101000100;
assign Simbolo[10][49] = 9'b100000000;
assign Simbolo[10][50] = 9'b100000000;
assign Simbolo[10][51] = 9'b100000000;
assign Simbolo[10][52] = 9'b100000000;
assign Simbolo[11][11] = 9'b100000000;
assign Simbolo[11][12] = 9'b101100100;
assign Simbolo[11][13] = 9'b111110001;
assign Simbolo[11][15] = 9'b100000000;
assign Simbolo[11][16] = 9'b100000000;
assign Simbolo[11][17] = 9'b100000000;
assign Simbolo[11][18] = 9'b100000000;
assign Simbolo[11][19] = 9'b100000000;
assign Simbolo[11][20] = 9'b100000000;
assign Simbolo[11][21] = 9'b101101000;
assign Simbolo[11][31] = 9'b100000000;
assign Simbolo[11][32] = 9'b100000000;
assign Simbolo[11][33] = 9'b100000000;
assign Simbolo[11][34] = 9'b100000000;
assign Simbolo[11][35] = 9'b100000000;
assign Simbolo[11][36] = 9'b100000000;
assign Simbolo[11][37] = 9'b100000000;
assign Simbolo[11][38] = 9'b100000000;
assign Simbolo[11][48] = 9'b101101000;
assign Simbolo[11][49] = 9'b100000000;
assign Simbolo[11][50] = 9'b100000000;
assign Simbolo[11][51] = 9'b100000000;
assign Simbolo[11][52] = 9'b100000000;
assign Simbolo[11][53] = 9'b100000000;
assign Simbolo[11][54] = 9'b100000000;
assign Simbolo[11][57] = 9'b101001000;
assign Simbolo[11][58] = 9'b100000000;
assign Simbolo[12][9] = 9'b100000000;
assign Simbolo[12][10] = 9'b100000000;
assign Simbolo[12][11] = 9'b100000000;
assign Simbolo[12][12] = 9'b101000100;
assign Simbolo[12][13] = 9'b101101000;
assign Simbolo[12][14] = 9'b100000000;
assign Simbolo[12][15] = 9'b100000000;
assign Simbolo[12][16] = 9'b100000000;
assign Simbolo[12][17] = 9'b100000000;
assign Simbolo[12][18] = 9'b100000000;
assign Simbolo[12][19] = 9'b100000000;
assign Simbolo[12][20] = 9'b100000000;
assign Simbolo[12][21] = 9'b100100100;
assign Simbolo[12][31] = 9'b100000000;
assign Simbolo[12][32] = 9'b100000000;
assign Simbolo[12][33] = 9'b100000000;
assign Simbolo[12][34] = 9'b101000000;
assign Simbolo[12][35] = 9'b100100000;
assign Simbolo[12][36] = 9'b100000000;
assign Simbolo[12][37] = 9'b100000000;
assign Simbolo[12][38] = 9'b100000000;
assign Simbolo[12][48] = 9'b100100100;
assign Simbolo[12][49] = 9'b100000000;
assign Simbolo[12][50] = 9'b100000000;
assign Simbolo[12][51] = 9'b100000000;
assign Simbolo[12][52] = 9'b100000000;
assign Simbolo[12][53] = 9'b100000000;
assign Simbolo[12][54] = 9'b100000000;
assign Simbolo[12][55] = 9'b100000000;
assign Simbolo[12][56] = 9'b101101000;
assign Simbolo[12][57] = 9'b101000100;
assign Simbolo[12][58] = 9'b100000000;
assign Simbolo[12][59] = 9'b100000000;
assign Simbolo[12][60] = 9'b100000000;
assign Simbolo[13][7] = 9'b100000000;
assign Simbolo[13][8] = 9'b100000000;
assign Simbolo[13][9] = 9'b100000000;
assign Simbolo[13][10] = 9'b100000000;
assign Simbolo[13][11] = 9'b100000000;
assign Simbolo[13][12] = 9'b100000000;
assign Simbolo[13][13] = 9'b101100100;
assign Simbolo[13][14] = 9'b100100000;
assign Simbolo[13][15] = 9'b100000000;
assign Simbolo[13][16] = 9'b100000000;
assign Simbolo[13][17] = 9'b100000000;
assign Simbolo[13][18] = 9'b100000000;
assign Simbolo[13][19] = 9'b100000000;
assign Simbolo[13][20] = 9'b100000000;
assign Simbolo[13][21] = 9'b100000000;
assign Simbolo[13][22] = 9'b100000000;
assign Simbolo[13][31] = 9'b100000000;
assign Simbolo[13][32] = 9'b100000000;
assign Simbolo[13][33] = 9'b100100000;
assign Simbolo[13][34] = 9'b101000000;
assign Simbolo[13][35] = 9'b101000000;
assign Simbolo[13][36] = 9'b100100000;
assign Simbolo[13][37] = 9'b100000000;
assign Simbolo[13][38] = 9'b100000000;
assign Simbolo[13][47] = 9'b100000000;
assign Simbolo[13][48] = 9'b100000000;
assign Simbolo[13][49] = 9'b100000000;
assign Simbolo[13][50] = 9'b100000000;
assign Simbolo[13][51] = 9'b100000000;
assign Simbolo[13][52] = 9'b100000000;
assign Simbolo[13][53] = 9'b100000000;
assign Simbolo[13][54] = 9'b100000000;
assign Simbolo[13][55] = 9'b100000000;
assign Simbolo[13][56] = 9'b101000100;
assign Simbolo[13][57] = 9'b100000000;
assign Simbolo[13][58] = 9'b100000000;
assign Simbolo[13][59] = 9'b100000000;
assign Simbolo[13][60] = 9'b100000000;
assign Simbolo[13][61] = 9'b100000000;
assign Simbolo[14][6] = 9'b100000000;
assign Simbolo[14][7] = 9'b100000000;
assign Simbolo[14][8] = 9'b100000000;
assign Simbolo[14][9] = 9'b100000000;
assign Simbolo[14][10] = 9'b100000000;
assign Simbolo[14][11] = 9'b100000000;
assign Simbolo[14][12] = 9'b100000000;
assign Simbolo[14][13] = 9'b100000000;
assign Simbolo[14][14] = 9'b101000000;
assign Simbolo[14][15] = 9'b100100000;
assign Simbolo[14][16] = 9'b100000000;
assign Simbolo[14][17] = 9'b100000000;
assign Simbolo[14][18] = 9'b100000000;
assign Simbolo[14][19] = 9'b100000000;
assign Simbolo[14][20] = 9'b100000000;
assign Simbolo[14][21] = 9'b100000000;
assign Simbolo[14][22] = 9'b100000000;
assign Simbolo[14][23] = 9'b100000000;
assign Simbolo[14][30] = 9'b100000000;
assign Simbolo[14][31] = 9'b100000000;
assign Simbolo[14][32] = 9'b100000000;
assign Simbolo[14][33] = 9'b101100000;
assign Simbolo[14][34] = 9'b100100000;
assign Simbolo[14][35] = 9'b100100000;
assign Simbolo[14][36] = 9'b101100000;
assign Simbolo[14][37] = 9'b100000000;
assign Simbolo[14][38] = 9'b100000000;
assign Simbolo[14][39] = 9'b100000000;
assign Simbolo[14][46] = 9'b100000000;
assign Simbolo[14][47] = 9'b100000000;
assign Simbolo[14][48] = 9'b100000000;
assign Simbolo[14][49] = 9'b100000000;
assign Simbolo[14][50] = 9'b100000000;
assign Simbolo[14][51] = 9'b100000000;
assign Simbolo[14][52] = 9'b100000000;
assign Simbolo[14][53] = 9'b100000000;
assign Simbolo[14][54] = 9'b100000000;
assign Simbolo[14][55] = 9'b100100000;
assign Simbolo[14][56] = 9'b100000000;
assign Simbolo[14][57] = 9'b100000000;
assign Simbolo[14][58] = 9'b100000000;
assign Simbolo[14][59] = 9'b100000000;
assign Simbolo[14][60] = 9'b100000000;
assign Simbolo[14][61] = 9'b100000000;
assign Simbolo[14][62] = 9'b100000000;
assign Simbolo[14][63] = 9'b100000000;
assign Simbolo[15][5] = 9'b100000000;
assign Simbolo[15][6] = 9'b100000000;
assign Simbolo[15][7] = 9'b100000000;
assign Simbolo[15][8] = 9'b100000000;
assign Simbolo[15][9] = 9'b100000000;
assign Simbolo[15][10] = 9'b100000000;
assign Simbolo[15][11] = 9'b100000000;
assign Simbolo[15][12] = 9'b100000000;
assign Simbolo[15][13] = 9'b100000000;
assign Simbolo[15][14] = 9'b100000000;
assign Simbolo[15][15] = 9'b100100000;
assign Simbolo[15][16] = 9'b100100000;
assign Simbolo[15][17] = 9'b100000000;
assign Simbolo[15][18] = 9'b100000000;
assign Simbolo[15][19] = 9'b100000000;
assign Simbolo[15][20] = 9'b100000000;
assign Simbolo[15][21] = 9'b100000000;
assign Simbolo[15][22] = 9'b100000000;
assign Simbolo[15][23] = 9'b100000000;
assign Simbolo[15][24] = 9'b100000000;
assign Simbolo[15][25] = 9'b100000000;
assign Simbolo[15][26] = 9'b100000000;
assign Simbolo[15][27] = 9'b100000000;
assign Simbolo[15][28] = 9'b100000000;
assign Simbolo[15][29] = 9'b100000000;
assign Simbolo[15][30] = 9'b100000000;
assign Simbolo[15][31] = 9'b100000000;
assign Simbolo[15][32] = 9'b101100000;
assign Simbolo[15][33] = 9'b101100100;
assign Simbolo[15][34] = 9'b100000000;
assign Simbolo[15][35] = 9'b100000000;
assign Simbolo[15][36] = 9'b101100100;
assign Simbolo[15][37] = 9'b101100000;
assign Simbolo[15][38] = 9'b100000000;
assign Simbolo[15][39] = 9'b100000000;
assign Simbolo[15][40] = 9'b100000000;
assign Simbolo[15][41] = 9'b100000000;
assign Simbolo[15][43] = 9'b100000000;
assign Simbolo[15][44] = 9'b100000000;
assign Simbolo[15][45] = 9'b100000000;
assign Simbolo[15][46] = 9'b100000000;
assign Simbolo[15][47] = 9'b100000000;
assign Simbolo[15][48] = 9'b100000000;
assign Simbolo[15][49] = 9'b100000000;
assign Simbolo[15][50] = 9'b100000000;
assign Simbolo[15][51] = 9'b100000000;
assign Simbolo[15][52] = 9'b100000000;
assign Simbolo[15][53] = 9'b100000000;
assign Simbolo[15][54] = 9'b100100000;
assign Simbolo[15][55] = 9'b100000000;
assign Simbolo[15][56] = 9'b100000000;
assign Simbolo[15][57] = 9'b100000000;
assign Simbolo[15][58] = 9'b100000000;
assign Simbolo[15][59] = 9'b100000000;
assign Simbolo[15][60] = 9'b100000000;
assign Simbolo[15][61] = 9'b100000000;
assign Simbolo[15][62] = 9'b100000000;
assign Simbolo[15][63] = 9'b100000000;
assign Simbolo[15][64] = 9'b100000000;
assign Simbolo[16][4] = 9'b100000000;
assign Simbolo[16][5] = 9'b100000000;
assign Simbolo[16][6] = 9'b100000000;
assign Simbolo[16][7] = 9'b100000000;
assign Simbolo[16][8] = 9'b100000000;
assign Simbolo[16][9] = 9'b100000000;
assign Simbolo[16][10] = 9'b100000000;
assign Simbolo[16][11] = 9'b100000000;
assign Simbolo[16][12] = 9'b100000000;
assign Simbolo[16][13] = 9'b100000000;
assign Simbolo[16][14] = 9'b100000000;
assign Simbolo[16][15] = 9'b100000000;
assign Simbolo[16][16] = 9'b100000000;
assign Simbolo[16][17] = 9'b100100000;
assign Simbolo[16][18] = 9'b100000000;
assign Simbolo[16][19] = 9'b100000000;
assign Simbolo[16][20] = 9'b100000000;
assign Simbolo[16][21] = 9'b100000000;
assign Simbolo[16][22] = 9'b100000000;
assign Simbolo[16][23] = 9'b100000000;
assign Simbolo[16][24] = 9'b100000000;
assign Simbolo[16][25] = 9'b100000000;
assign Simbolo[16][26] = 9'b100000000;
assign Simbolo[16][27] = 9'b100000000;
assign Simbolo[16][28] = 9'b100000000;
assign Simbolo[16][29] = 9'b100000000;
assign Simbolo[16][30] = 9'b100000000;
assign Simbolo[16][31] = 9'b101100000;
assign Simbolo[16][32] = 9'b111101000;
assign Simbolo[16][33] = 9'b100100100;
assign Simbolo[16][34] = 9'b100000000;
assign Simbolo[16][35] = 9'b100000000;
assign Simbolo[16][36] = 9'b101000100;
assign Simbolo[16][37] = 9'b111101000;
assign Simbolo[16][38] = 9'b101000000;
assign Simbolo[16][39] = 9'b100000000;
assign Simbolo[16][40] = 9'b100000000;
assign Simbolo[16][41] = 9'b100000000;
assign Simbolo[16][42] = 9'b100000000;
assign Simbolo[16][43] = 9'b100000000;
assign Simbolo[16][44] = 9'b100000000;
assign Simbolo[16][45] = 9'b100000000;
assign Simbolo[16][46] = 9'b100000000;
assign Simbolo[16][47] = 9'b100000000;
assign Simbolo[16][48] = 9'b100000000;
assign Simbolo[16][49] = 9'b100000000;
assign Simbolo[16][50] = 9'b100000000;
assign Simbolo[16][51] = 9'b100000000;
assign Simbolo[16][52] = 9'b100000000;
assign Simbolo[16][53] = 9'b100000000;
assign Simbolo[16][54] = 9'b100000000;
assign Simbolo[16][55] = 9'b100000000;
assign Simbolo[16][56] = 9'b100000000;
assign Simbolo[16][57] = 9'b100000000;
assign Simbolo[16][58] = 9'b100000000;
assign Simbolo[16][59] = 9'b100000000;
assign Simbolo[16][60] = 9'b100000000;
assign Simbolo[16][61] = 9'b100000000;
assign Simbolo[16][62] = 9'b100000000;
assign Simbolo[16][63] = 9'b100000000;
assign Simbolo[16][64] = 9'b100000000;
assign Simbolo[16][65] = 9'b100000000;
assign Simbolo[17][3] = 9'b100000000;
assign Simbolo[17][4] = 9'b100000000;
assign Simbolo[17][5] = 9'b100000000;
assign Simbolo[17][6] = 9'b100000000;
assign Simbolo[17][7] = 9'b100000000;
assign Simbolo[17][8] = 9'b100000000;
assign Simbolo[17][9] = 9'b100000000;
assign Simbolo[17][10] = 9'b100000000;
assign Simbolo[17][11] = 9'b100000000;
assign Simbolo[17][12] = 9'b100000000;
assign Simbolo[17][13] = 9'b100000000;
assign Simbolo[17][14] = 9'b100000000;
assign Simbolo[17][15] = 9'b100000000;
assign Simbolo[17][16] = 9'b100000000;
assign Simbolo[17][17] = 9'b100000000;
assign Simbolo[17][18] = 9'b100000000;
assign Simbolo[17][19] = 9'b100000000;
assign Simbolo[17][20] = 9'b100000000;
assign Simbolo[17][21] = 9'b100000000;
assign Simbolo[17][22] = 9'b100000000;
assign Simbolo[17][23] = 9'b100000000;
assign Simbolo[17][24] = 9'b100000000;
assign Simbolo[17][25] = 9'b100000000;
assign Simbolo[17][26] = 9'b100000000;
assign Simbolo[17][27] = 9'b100000000;
assign Simbolo[17][28] = 9'b100000000;
assign Simbolo[17][29] = 9'b100100000;
assign Simbolo[17][30] = 9'b101100100;
assign Simbolo[17][31] = 9'b111101000;
assign Simbolo[17][32] = 9'b110001000;
assign Simbolo[17][33] = 9'b100000000;
assign Simbolo[17][34] = 9'b100000000;
assign Simbolo[17][35] = 9'b100000000;
assign Simbolo[17][36] = 9'b100000000;
assign Simbolo[17][37] = 9'b110001000;
assign Simbolo[17][38] = 9'b111101000;
assign Simbolo[17][39] = 9'b101100000;
assign Simbolo[17][40] = 9'b100100000;
assign Simbolo[17][41] = 9'b100000000;
assign Simbolo[17][42] = 9'b100000000;
assign Simbolo[17][43] = 9'b100000000;
assign Simbolo[17][44] = 9'b100000000;
assign Simbolo[17][45] = 9'b100000000;
assign Simbolo[17][46] = 9'b100000000;
assign Simbolo[17][47] = 9'b100000000;
assign Simbolo[17][48] = 9'b100000000;
assign Simbolo[17][49] = 9'b100000000;
assign Simbolo[17][50] = 9'b100000000;
assign Simbolo[17][51] = 9'b100000000;
assign Simbolo[17][52] = 9'b100000000;
assign Simbolo[17][53] = 9'b100000000;
assign Simbolo[17][54] = 9'b100000000;
assign Simbolo[17][55] = 9'b100000000;
assign Simbolo[17][56] = 9'b100000000;
assign Simbolo[17][57] = 9'b100000000;
assign Simbolo[17][58] = 9'b100000000;
assign Simbolo[17][59] = 9'b100000000;
assign Simbolo[17][60] = 9'b100000000;
assign Simbolo[17][61] = 9'b100000000;
assign Simbolo[17][62] = 9'b100000000;
assign Simbolo[17][63] = 9'b100000000;
assign Simbolo[17][64] = 9'b100000000;
assign Simbolo[17][65] = 9'b100000000;
assign Simbolo[17][66] = 9'b100000000;
assign Simbolo[18][3] = 9'b100000000;
assign Simbolo[18][4] = 9'b100000000;
assign Simbolo[18][5] = 9'b100000000;
assign Simbolo[18][6] = 9'b100000000;
assign Simbolo[18][7] = 9'b100000000;
assign Simbolo[18][8] = 9'b100000000;
assign Simbolo[18][9] = 9'b100000000;
assign Simbolo[18][10] = 9'b100000000;
assign Simbolo[18][11] = 9'b100000000;
assign Simbolo[18][12] = 9'b100000000;
assign Simbolo[18][13] = 9'b100000000;
assign Simbolo[18][14] = 9'b100000000;
assign Simbolo[18][15] = 9'b100000000;
assign Simbolo[18][16] = 9'b100000000;
assign Simbolo[18][17] = 9'b100000000;
assign Simbolo[18][18] = 9'b100000000;
assign Simbolo[18][19] = 9'b100000000;
assign Simbolo[18][20] = 9'b100000000;
assign Simbolo[18][21] = 9'b100000000;
assign Simbolo[18][22] = 9'b100000000;
assign Simbolo[18][23] = 9'b100000000;
assign Simbolo[18][24] = 9'b100000000;
assign Simbolo[18][25] = 9'b100000000;
assign Simbolo[18][26] = 9'b100100000;
assign Simbolo[18][27] = 9'b100100000;
assign Simbolo[18][28] = 9'b101000000;
assign Simbolo[18][29] = 9'b110000100;
assign Simbolo[18][30] = 9'b110101000;
assign Simbolo[18][31] = 9'b101101000;
assign Simbolo[18][32] = 9'b100000000;
assign Simbolo[18][33] = 9'b100000000;
assign Simbolo[18][34] = 9'b100000000;
assign Simbolo[18][35] = 9'b100000000;
assign Simbolo[18][36] = 9'b100000000;
assign Simbolo[18][37] = 9'b100000000;
assign Simbolo[18][38] = 9'b110001000;
assign Simbolo[18][39] = 9'b110101000;
assign Simbolo[18][40] = 9'b110000100;
assign Simbolo[18][41] = 9'b101000000;
assign Simbolo[18][42] = 9'b100100000;
assign Simbolo[18][43] = 9'b100000000;
assign Simbolo[18][44] = 9'b100000000;
assign Simbolo[18][45] = 9'b100000000;
assign Simbolo[18][46] = 9'b100000000;
assign Simbolo[18][47] = 9'b100000000;
assign Simbolo[18][48] = 9'b100000000;
assign Simbolo[18][49] = 9'b100000000;
assign Simbolo[18][50] = 9'b100000000;
assign Simbolo[18][51] = 9'b100000000;
assign Simbolo[18][52] = 9'b100000000;
assign Simbolo[18][53] = 9'b100000000;
assign Simbolo[18][54] = 9'b100000000;
assign Simbolo[18][55] = 9'b100000000;
assign Simbolo[18][56] = 9'b100000000;
assign Simbolo[18][57] = 9'b100000000;
assign Simbolo[18][58] = 9'b100000000;
assign Simbolo[18][59] = 9'b100000000;
assign Simbolo[18][60] = 9'b100000000;
assign Simbolo[18][61] = 9'b100000000;
assign Simbolo[18][62] = 9'b100000000;
assign Simbolo[18][63] = 9'b100000000;
assign Simbolo[18][64] = 9'b100000000;
assign Simbolo[18][65] = 9'b100000000;
assign Simbolo[18][66] = 9'b100000000;
assign Simbolo[19][2] = 9'b100000000;
assign Simbolo[19][3] = 9'b100000000;
assign Simbolo[19][4] = 9'b100000000;
assign Simbolo[19][5] = 9'b100000000;
assign Simbolo[19][6] = 9'b100000000;
assign Simbolo[19][7] = 9'b100000000;
assign Simbolo[19][8] = 9'b100000000;
assign Simbolo[19][9] = 9'b100000000;
assign Simbolo[19][10] = 9'b100000000;
assign Simbolo[19][11] = 9'b100100000;
assign Simbolo[19][12] = 9'b100100000;
assign Simbolo[19][13] = 9'b100100000;
assign Simbolo[19][14] = 9'b100000000;
assign Simbolo[19][15] = 9'b100000000;
assign Simbolo[19][16] = 9'b100000000;
assign Simbolo[19][17] = 9'b100000000;
assign Simbolo[19][18] = 9'b100000000;
assign Simbolo[19][19] = 9'b100000000;
assign Simbolo[19][20] = 9'b100000000;
assign Simbolo[19][21] = 9'b100000000;
assign Simbolo[19][22] = 9'b100000000;
assign Simbolo[19][23] = 9'b100000000;
assign Simbolo[19][24] = 9'b100000000;
assign Simbolo[19][25] = 9'b100000000;
assign Simbolo[19][26] = 9'b100000000;
assign Simbolo[19][27] = 9'b100000000;
assign Simbolo[19][28] = 9'b100000000;
assign Simbolo[19][29] = 9'b100000000;
assign Simbolo[19][30] = 9'b100000000;
assign Simbolo[19][31] = 9'b100000000;
assign Simbolo[19][32] = 9'b100000000;
assign Simbolo[19][33] = 9'b100000000;
assign Simbolo[19][34] = 9'b100000000;
assign Simbolo[19][35] = 9'b100000000;
assign Simbolo[19][36] = 9'b100000000;
assign Simbolo[19][37] = 9'b100000000;
assign Simbolo[19][38] = 9'b100000000;
assign Simbolo[19][39] = 9'b100000000;
assign Simbolo[19][40] = 9'b100100000;
assign Simbolo[19][41] = 9'b100100000;
assign Simbolo[19][42] = 9'b100000000;
assign Simbolo[19][43] = 9'b100000000;
assign Simbolo[19][44] = 9'b100000000;
assign Simbolo[19][45] = 9'b100000000;
assign Simbolo[19][46] = 9'b100000000;
assign Simbolo[19][47] = 9'b100000000;
assign Simbolo[19][48] = 9'b100000000;
assign Simbolo[19][49] = 9'b100000000;
assign Simbolo[19][50] = 9'b100000000;
assign Simbolo[19][51] = 9'b100000000;
assign Simbolo[19][52] = 9'b100000000;
assign Simbolo[19][53] = 9'b100000000;
assign Simbolo[19][54] = 9'b100000000;
assign Simbolo[19][55] = 9'b100000000;
assign Simbolo[19][56] = 9'b100000000;
assign Simbolo[19][57] = 9'b100000000;
assign Simbolo[19][58] = 9'b100000000;
assign Simbolo[19][59] = 9'b100000000;
assign Simbolo[19][60] = 9'b100000000;
assign Simbolo[19][61] = 9'b100000000;
assign Simbolo[19][62] = 9'b100000000;
assign Simbolo[19][63] = 9'b100000000;
assign Simbolo[19][64] = 9'b100000000;
assign Simbolo[19][65] = 9'b100000000;
assign Simbolo[19][66] = 9'b100000000;
assign Simbolo[19][67] = 9'b100000000;
assign Simbolo[20][2] = 9'b100000000;
assign Simbolo[20][3] = 9'b100000000;
assign Simbolo[20][4] = 9'b100000000;
assign Simbolo[20][5] = 9'b100000000;
assign Simbolo[20][6] = 9'b100000000;
assign Simbolo[20][7] = 9'b100000000;
assign Simbolo[20][8] = 9'b100000000;
assign Simbolo[20][9] = 9'b100100000;
assign Simbolo[20][10] = 9'b101000000;
assign Simbolo[20][11] = 9'b100100000;
assign Simbolo[20][12] = 9'b100000000;
assign Simbolo[20][13] = 9'b100000000;
assign Simbolo[20][14] = 9'b100000000;
assign Simbolo[20][15] = 9'b100000000;
assign Simbolo[20][16] = 9'b100000000;
assign Simbolo[20][17] = 9'b100000000;
assign Simbolo[20][18] = 9'b100000000;
assign Simbolo[20][19] = 9'b100000000;
assign Simbolo[20][20] = 9'b100000000;
assign Simbolo[20][21] = 9'b100000000;
assign Simbolo[20][22] = 9'b100000000;
assign Simbolo[20][23] = 9'b100000000;
assign Simbolo[20][24] = 9'b100000000;
assign Simbolo[20][25] = 9'b100000000;
assign Simbolo[20][26] = 9'b100000000;
assign Simbolo[20][27] = 9'b100000000;
assign Simbolo[20][28] = 9'b100000000;
assign Simbolo[20][29] = 9'b100000000;
assign Simbolo[20][30] = 9'b100000000;
assign Simbolo[20][31] = 9'b100000000;
assign Simbolo[20][32] = 9'b100000000;
assign Simbolo[20][33] = 9'b100000000;
assign Simbolo[20][34] = 9'b100000000;
assign Simbolo[20][35] = 9'b100000000;
assign Simbolo[20][36] = 9'b100000000;
assign Simbolo[20][37] = 9'b100000000;
assign Simbolo[20][38] = 9'b100000000;
assign Simbolo[20][39] = 9'b100000000;
assign Simbolo[20][40] = 9'b100000000;
assign Simbolo[20][41] = 9'b100000000;
assign Simbolo[20][42] = 9'b100000000;
assign Simbolo[20][43] = 9'b100000000;
assign Simbolo[20][44] = 9'b100000000;
assign Simbolo[20][45] = 9'b100000000;
assign Simbolo[20][46] = 9'b100000000;
assign Simbolo[20][47] = 9'b100000000;
assign Simbolo[20][48] = 9'b100000000;
assign Simbolo[20][49] = 9'b100000000;
assign Simbolo[20][50] = 9'b100000000;
assign Simbolo[20][51] = 9'b100000000;
assign Simbolo[20][52] = 9'b100000000;
assign Simbolo[20][53] = 9'b100000000;
assign Simbolo[20][54] = 9'b100000000;
assign Simbolo[20][55] = 9'b100000000;
assign Simbolo[20][56] = 9'b100000000;
assign Simbolo[20][57] = 9'b100000000;
assign Simbolo[20][58] = 9'b100100000;
assign Simbolo[20][59] = 9'b101000000;
assign Simbolo[20][60] = 9'b100000000;
assign Simbolo[20][61] = 9'b100000000;
assign Simbolo[20][62] = 9'b100000000;
assign Simbolo[20][63] = 9'b100000000;
assign Simbolo[20][64] = 9'b100000000;
assign Simbolo[20][65] = 9'b100000000;
assign Simbolo[20][66] = 9'b100000000;
assign Simbolo[20][67] = 9'b100000000;
assign Simbolo[21][2] = 9'b100000000;
assign Simbolo[21][3] = 9'b100000000;
assign Simbolo[21][4] = 9'b100000000;
assign Simbolo[21][5] = 9'b100000000;
assign Simbolo[21][6] = 9'b100000000;
assign Simbolo[21][7] = 9'b100000000;
assign Simbolo[21][8] = 9'b101000000;
assign Simbolo[21][9] = 9'b101000000;
assign Simbolo[21][10] = 9'b100000000;
assign Simbolo[21][11] = 9'b100000000;
assign Simbolo[21][12] = 9'b100000000;
assign Simbolo[21][13] = 9'b100000000;
assign Simbolo[21][14] = 9'b100000000;
assign Simbolo[21][15] = 9'b100000000;
assign Simbolo[21][16] = 9'b100000000;
assign Simbolo[21][17] = 9'b100000000;
assign Simbolo[21][18] = 9'b100000000;
assign Simbolo[21][19] = 9'b100000000;
assign Simbolo[21][20] = 9'b100000000;
assign Simbolo[21][21] = 9'b100000000;
assign Simbolo[21][22] = 9'b100000000;
assign Simbolo[21][23] = 9'b100000000;
assign Simbolo[21][24] = 9'b100000000;
assign Simbolo[21][25] = 9'b100000000;
assign Simbolo[21][26] = 9'b100000000;
assign Simbolo[21][27] = 9'b100000000;
assign Simbolo[21][28] = 9'b100000000;
assign Simbolo[21][29] = 9'b100000000;
assign Simbolo[21][30] = 9'b100000000;
assign Simbolo[21][31] = 9'b100000000;
assign Simbolo[21][32] = 9'b100000000;
assign Simbolo[21][33] = 9'b100000000;
assign Simbolo[21][34] = 9'b100000000;
assign Simbolo[21][35] = 9'b100000000;
assign Simbolo[21][36] = 9'b100000000;
assign Simbolo[21][37] = 9'b100000000;
assign Simbolo[21][38] = 9'b100000000;
assign Simbolo[21][39] = 9'b100000000;
assign Simbolo[21][40] = 9'b100000000;
assign Simbolo[21][41] = 9'b100000000;
assign Simbolo[21][42] = 9'b100000000;
assign Simbolo[21][43] = 9'b100000000;
assign Simbolo[21][44] = 9'b100000000;
assign Simbolo[21][45] = 9'b100000000;
assign Simbolo[21][46] = 9'b100000000;
assign Simbolo[21][47] = 9'b100000000;
assign Simbolo[21][48] = 9'b100000000;
assign Simbolo[21][49] = 9'b100000000;
assign Simbolo[21][50] = 9'b100000000;
assign Simbolo[21][51] = 9'b100000000;
assign Simbolo[21][52] = 9'b100000000;
assign Simbolo[21][53] = 9'b100000000;
assign Simbolo[21][54] = 9'b100000000;
assign Simbolo[21][55] = 9'b100000000;
assign Simbolo[21][56] = 9'b100000000;
assign Simbolo[21][57] = 9'b100000000;
assign Simbolo[21][58] = 9'b100000000;
assign Simbolo[21][59] = 9'b100000000;
assign Simbolo[21][60] = 9'b101000000;
assign Simbolo[21][61] = 9'b100100000;
assign Simbolo[21][62] = 9'b100000000;
assign Simbolo[21][63] = 9'b100000000;
assign Simbolo[21][64] = 9'b100000000;
assign Simbolo[21][65] = 9'b100000000;
assign Simbolo[21][66] = 9'b100000000;
assign Simbolo[21][67] = 9'b100000000;
assign Simbolo[22][2] = 9'b100000000;
assign Simbolo[22][3] = 9'b100000000;
assign Simbolo[22][4] = 9'b100000000;
assign Simbolo[22][5] = 9'b100000000;
assign Simbolo[22][6] = 9'b100000000;
assign Simbolo[22][7] = 9'b100100000;
assign Simbolo[22][8] = 9'b101100100;
assign Simbolo[22][9] = 9'b100000000;
assign Simbolo[22][10] = 9'b100000000;
assign Simbolo[22][11] = 9'b100000000;
assign Simbolo[22][12] = 9'b100000000;
assign Simbolo[22][13] = 9'b100000000;
assign Simbolo[22][14] = 9'b100000000;
assign Simbolo[22][15] = 9'b100000000;
assign Simbolo[22][16] = 9'b100000000;
assign Simbolo[22][17] = 9'b100000000;
assign Simbolo[22][18] = 9'b100000000;
assign Simbolo[22][19] = 9'b100000000;
assign Simbolo[22][20] = 9'b100000000;
assign Simbolo[22][21] = 9'b100000000;
assign Simbolo[22][22] = 9'b100000000;
assign Simbolo[22][23] = 9'b100000000;
assign Simbolo[22][24] = 9'b100000000;
assign Simbolo[22][25] = 9'b100000000;
assign Simbolo[22][26] = 9'b100000000;
assign Simbolo[22][27] = 9'b100000000;
assign Simbolo[22][28] = 9'b100100000;
assign Simbolo[22][29] = 9'b100100000;
assign Simbolo[22][30] = 9'b100000000;
assign Simbolo[22][31] = 9'b100000000;
assign Simbolo[22][32] = 9'b100000000;
assign Simbolo[22][33] = 9'b100000000;
assign Simbolo[22][34] = 9'b100000000;
assign Simbolo[22][35] = 9'b100000000;
assign Simbolo[22][36] = 9'b100000000;
assign Simbolo[22][37] = 9'b100000000;
assign Simbolo[22][38] = 9'b100000000;
assign Simbolo[22][39] = 9'b100000000;
assign Simbolo[22][40] = 9'b100100000;
assign Simbolo[22][41] = 9'b100100000;
assign Simbolo[22][42] = 9'b100000000;
assign Simbolo[22][43] = 9'b100000000;
assign Simbolo[22][44] = 9'b100000000;
assign Simbolo[22][45] = 9'b100000000;
assign Simbolo[22][46] = 9'b100000000;
assign Simbolo[22][47] = 9'b100000000;
assign Simbolo[22][48] = 9'b100000000;
assign Simbolo[22][49] = 9'b100000000;
assign Simbolo[22][50] = 9'b100000000;
assign Simbolo[22][51] = 9'b100000000;
assign Simbolo[22][52] = 9'b100000000;
assign Simbolo[22][53] = 9'b100000000;
assign Simbolo[22][54] = 9'b100000000;
assign Simbolo[22][55] = 9'b100000000;
assign Simbolo[22][56] = 9'b100000000;
assign Simbolo[22][57] = 9'b100000000;
assign Simbolo[22][58] = 9'b100000000;
assign Simbolo[22][59] = 9'b100000000;
assign Simbolo[22][60] = 9'b100000000;
assign Simbolo[22][61] = 9'b101100100;
assign Simbolo[22][62] = 9'b100100000;
assign Simbolo[22][63] = 9'b100000000;
assign Simbolo[22][64] = 9'b100000000;
assign Simbolo[22][65] = 9'b100000000;
assign Simbolo[22][66] = 9'b100000000;
assign Simbolo[22][67] = 9'b100000000;
assign Simbolo[23][3] = 9'b100000000;
assign Simbolo[23][4] = 9'b100000000;
assign Simbolo[23][5] = 9'b100000000;
assign Simbolo[23][6] = 9'b100000000;
assign Simbolo[23][7] = 9'b101100100;
assign Simbolo[23][8] = 9'b101000100;
assign Simbolo[23][9] = 9'b100000000;
assign Simbolo[23][10] = 9'b100000000;
assign Simbolo[23][11] = 9'b100000000;
assign Simbolo[23][12] = 9'b100000000;
assign Simbolo[23][13] = 9'b100000000;
assign Simbolo[23][14] = 9'b100000000;
assign Simbolo[23][15] = 9'b100000000;
assign Simbolo[23][16] = 9'b100000000;
assign Simbolo[23][17] = 9'b100000000;
assign Simbolo[23][18] = 9'b100000000;
assign Simbolo[23][19] = 9'b100000000;
assign Simbolo[23][20] = 9'b100000000;
assign Simbolo[23][21] = 9'b100000000;
assign Simbolo[23][22] = 9'b100000000;
assign Simbolo[23][23] = 9'b100000000;
assign Simbolo[23][24] = 9'b100000000;
assign Simbolo[23][25] = 9'b100000000;
assign Simbolo[23][26] = 9'b100000000;
assign Simbolo[23][27] = 9'b100000000;
assign Simbolo[23][28] = 9'b100000000;
assign Simbolo[23][29] = 9'b101000000;
assign Simbolo[23][30] = 9'b101000000;
assign Simbolo[23][31] = 9'b100000000;
assign Simbolo[23][32] = 9'b100000000;
assign Simbolo[23][33] = 9'b100000000;
assign Simbolo[23][34] = 9'b100000000;
assign Simbolo[23][35] = 9'b100000000;
assign Simbolo[23][36] = 9'b100000000;
assign Simbolo[23][37] = 9'b100000000;
assign Simbolo[23][38] = 9'b100000000;
assign Simbolo[23][39] = 9'b101100000;
assign Simbolo[23][40] = 9'b101000000;
assign Simbolo[23][41] = 9'b100000000;
assign Simbolo[23][42] = 9'b100000000;
assign Simbolo[23][43] = 9'b100000000;
assign Simbolo[23][44] = 9'b100000000;
assign Simbolo[23][45] = 9'b100000000;
assign Simbolo[23][46] = 9'b100000000;
assign Simbolo[23][47] = 9'b100000000;
assign Simbolo[23][48] = 9'b100000000;
assign Simbolo[23][49] = 9'b100000000;
assign Simbolo[23][50] = 9'b100000000;
assign Simbolo[23][51] = 9'b100000000;
assign Simbolo[23][52] = 9'b100000000;
assign Simbolo[23][53] = 9'b100000000;
assign Simbolo[23][54] = 9'b100000000;
assign Simbolo[23][55] = 9'b100000000;
assign Simbolo[23][56] = 9'b100000000;
assign Simbolo[23][57] = 9'b100000000;
assign Simbolo[23][58] = 9'b100000000;
assign Simbolo[23][59] = 9'b100000000;
assign Simbolo[23][60] = 9'b100000000;
assign Simbolo[23][61] = 9'b101000100;
assign Simbolo[23][62] = 9'b101100100;
assign Simbolo[23][63] = 9'b100000000;
assign Simbolo[23][64] = 9'b100000000;
assign Simbolo[23][65] = 9'b100000000;
assign Simbolo[23][66] = 9'b100000000;
assign Simbolo[24][3] = 9'b100000000;
assign Simbolo[24][4] = 9'b100000000;
assign Simbolo[24][5] = 9'b100000000;
assign Simbolo[24][6] = 9'b100000000;
assign Simbolo[24][7] = 9'b110001000;
assign Simbolo[24][9] = 9'b100000000;
assign Simbolo[24][10] = 9'b100000000;
assign Simbolo[24][11] = 9'b100000000;
assign Simbolo[24][12] = 9'b100000000;
assign Simbolo[24][13] = 9'b100000000;
assign Simbolo[24][14] = 9'b100000000;
assign Simbolo[24][15] = 9'b100000000;
assign Simbolo[24][16] = 9'b100000000;
assign Simbolo[24][17] = 9'b100000000;
assign Simbolo[24][18] = 9'b100000000;
assign Simbolo[24][19] = 9'b100000000;
assign Simbolo[24][20] = 9'b100000000;
assign Simbolo[24][21] = 9'b100000000;
assign Simbolo[24][22] = 9'b100000000;
assign Simbolo[24][23] = 9'b100000000;
assign Simbolo[24][24] = 9'b100000000;
assign Simbolo[24][25] = 9'b100000000;
assign Simbolo[24][26] = 9'b100000000;
assign Simbolo[24][27] = 9'b100000000;
assign Simbolo[24][28] = 9'b100000000;
assign Simbolo[24][29] = 9'b100000000;
assign Simbolo[24][30] = 9'b101000000;
assign Simbolo[24][31] = 9'b110000100;
assign Simbolo[24][32] = 9'b100100000;
assign Simbolo[24][33] = 9'b100000000;
assign Simbolo[24][34] = 9'b100000000;
assign Simbolo[24][35] = 9'b100000000;
assign Simbolo[24][36] = 9'b100000000;
assign Simbolo[24][37] = 9'b101000000;
assign Simbolo[24][38] = 9'b110000100;
assign Simbolo[24][39] = 9'b101000000;
assign Simbolo[24][40] = 9'b100000000;
assign Simbolo[24][41] = 9'b100000000;
assign Simbolo[24][42] = 9'b100000000;
assign Simbolo[24][43] = 9'b100000000;
assign Simbolo[24][44] = 9'b100000000;
assign Simbolo[24][45] = 9'b100000000;
assign Simbolo[24][46] = 9'b100000000;
assign Simbolo[24][47] = 9'b100000000;
assign Simbolo[24][48] = 9'b100000000;
assign Simbolo[24][49] = 9'b100000000;
assign Simbolo[24][50] = 9'b100000000;
assign Simbolo[24][51] = 9'b100000000;
assign Simbolo[24][52] = 9'b100000000;
assign Simbolo[24][53] = 9'b100000000;
assign Simbolo[24][54] = 9'b100000000;
assign Simbolo[24][55] = 9'b100000000;
assign Simbolo[24][56] = 9'b100000000;
assign Simbolo[24][57] = 9'b100000000;
assign Simbolo[24][58] = 9'b100000000;
assign Simbolo[24][59] = 9'b100000000;
assign Simbolo[24][60] = 9'b100000000;
assign Simbolo[24][62] = 9'b101101000;
assign Simbolo[24][63] = 9'b100000000;
assign Simbolo[24][64] = 9'b100000000;
assign Simbolo[24][65] = 9'b100000000;
assign Simbolo[24][66] = 9'b100000000;
assign Simbolo[25][3] = 9'b100000000;
assign Simbolo[25][4] = 9'b100000000;
assign Simbolo[25][5] = 9'b100000000;
assign Simbolo[25][6] = 9'b100000000;
assign Simbolo[25][7] = 9'b101101000;
assign Simbolo[25][10] = 9'b100000000;
assign Simbolo[25][11] = 9'b100000000;
assign Simbolo[25][12] = 9'b100000000;
assign Simbolo[25][13] = 9'b100000000;
assign Simbolo[25][14] = 9'b100000000;
assign Simbolo[25][15] = 9'b100000000;
assign Simbolo[25][16] = 9'b100000000;
assign Simbolo[25][17] = 9'b100000000;
assign Simbolo[25][18] = 9'b100000000;
assign Simbolo[25][19] = 9'b100000000;
assign Simbolo[25][22] = 9'b100000000;
assign Simbolo[25][23] = 9'b100000000;
assign Simbolo[25][24] = 9'b100000000;
assign Simbolo[25][25] = 9'b100000000;
assign Simbolo[25][26] = 9'b100000000;
assign Simbolo[25][27] = 9'b100000000;
assign Simbolo[25][28] = 9'b100100000;
assign Simbolo[25][29] = 9'b100000000;
assign Simbolo[25][30] = 9'b100000000;
assign Simbolo[25][31] = 9'b101000000;
assign Simbolo[25][32] = 9'b110000100;
assign Simbolo[25][33] = 9'b101000000;
assign Simbolo[25][34] = 9'b100000000;
assign Simbolo[25][35] = 9'b100000000;
assign Simbolo[25][36] = 9'b101000100;
assign Simbolo[25][37] = 9'b110000100;
assign Simbolo[25][38] = 9'b101000000;
assign Simbolo[25][39] = 9'b100000000;
assign Simbolo[25][40] = 9'b100000000;
assign Simbolo[25][41] = 9'b100000000;
assign Simbolo[25][42] = 9'b100000000;
assign Simbolo[25][43] = 9'b100000000;
assign Simbolo[25][44] = 9'b100000000;
assign Simbolo[25][45] = 9'b100000000;
assign Simbolo[25][46] = 9'b100000000;
assign Simbolo[25][47] = 9'b100000000;
assign Simbolo[25][48] = 9'b100000000;
assign Simbolo[25][49] = 9'b100000000;
assign Simbolo[25][50] = 9'b100000000;
assign Simbolo[25][51] = 9'b100000000;
assign Simbolo[25][52] = 9'b100000000;
assign Simbolo[25][53] = 9'b100000000;
assign Simbolo[25][54] = 9'b100000000;
assign Simbolo[25][55] = 9'b100000000;
assign Simbolo[25][56] = 9'b100000000;
assign Simbolo[25][57] = 9'b100000000;
assign Simbolo[25][58] = 9'b100000000;
assign Simbolo[25][59] = 9'b100000000;
assign Simbolo[25][62] = 9'b101101000;
assign Simbolo[25][63] = 9'b100000000;
assign Simbolo[25][64] = 9'b100000000;
assign Simbolo[25][65] = 9'b100000000;
assign Simbolo[25][66] = 9'b100000000;
assign Simbolo[26][4] = 9'b100000000;
assign Simbolo[26][5] = 9'b100000000;
assign Simbolo[26][6] = 9'b100000000;
assign Simbolo[26][7] = 9'b101000100;
assign Simbolo[26][11] = 9'b100000000;
assign Simbolo[26][12] = 9'b100000000;
assign Simbolo[26][13] = 9'b100000000;
assign Simbolo[26][14] = 9'b100000000;
assign Simbolo[26][15] = 9'b100000000;
assign Simbolo[26][16] = 9'b100000000;
assign Simbolo[26][17] = 9'b101000100;
assign Simbolo[26][24] = 9'b100000000;
assign Simbolo[26][25] = 9'b100000000;
assign Simbolo[26][31] = 9'b100100000;
assign Simbolo[26][32] = 9'b101000000;
assign Simbolo[26][33] = 9'b110000100;
assign Simbolo[26][34] = 9'b100100000;
assign Simbolo[26][35] = 9'b100100000;
assign Simbolo[26][36] = 9'b110000100;
assign Simbolo[26][37] = 9'b100100000;
assign Simbolo[26][38] = 9'b100000000;
assign Simbolo[26][43] = 9'b100100100;
assign Simbolo[26][44] = 9'b100000000;
assign Simbolo[26][45] = 9'b100000000;
assign Simbolo[26][52] = 9'b100100000;
assign Simbolo[26][53] = 9'b100000000;
assign Simbolo[26][54] = 9'b100000000;
assign Simbolo[26][55] = 9'b100000000;
assign Simbolo[26][56] = 9'b100000000;
assign Simbolo[26][57] = 9'b100000000;
assign Simbolo[26][58] = 9'b100000000;
assign Simbolo[26][59] = 9'b100000000;
assign Simbolo[26][62] = 9'b101000100;
assign Simbolo[26][63] = 9'b100000000;
assign Simbolo[26][64] = 9'b100000000;
assign Simbolo[26][65] = 9'b100000000;
assign Simbolo[27][5] = 9'b100000000;
assign Simbolo[27][6] = 9'b100000000;
assign Simbolo[27][7] = 9'b100000000;
assign Simbolo[27][8] = 9'b110000100;
assign Simbolo[27][12] = 9'b100000000;
assign Simbolo[27][13] = 9'b100000000;
assign Simbolo[27][14] = 9'b100000000;
assign Simbolo[27][15] = 9'b100000000;
assign Simbolo[27][16] = 9'b100100000;
assign Simbolo[27][17] = 9'b110110001;
assign Simbolo[27][32] = 9'b100100000;
assign Simbolo[27][33] = 9'b101100000;
assign Simbolo[27][34] = 9'b101000000;
assign Simbolo[27][35] = 9'b101000000;
assign Simbolo[27][36] = 9'b101000000;
assign Simbolo[27][37] = 9'b100000000;
assign Simbolo[27][52] = 9'b110001101;
assign Simbolo[27][53] = 9'b100000000;
assign Simbolo[27][54] = 9'b100000000;
assign Simbolo[27][55] = 9'b100000000;
assign Simbolo[27][56] = 9'b100000000;
assign Simbolo[27][57] = 9'b100000000;
assign Simbolo[27][61] = 9'b101100100;
assign Simbolo[27][62] = 9'b100000000;
assign Simbolo[27][63] = 9'b100000000;
assign Simbolo[27][64] = 9'b100000000;
assign Simbolo[28][6] = 9'b100000000;
assign Simbolo[28][7] = 9'b100000000;
assign Simbolo[28][8] = 9'b100100000;
assign Simbolo[28][14] = 9'b100000000;
assign Simbolo[28][15] = 9'b100000000;
assign Simbolo[28][16] = 9'b100000000;
assign Simbolo[28][17] = 9'b101101001;
assign Simbolo[28][33] = 9'b101000000;
assign Simbolo[28][34] = 9'b101000000;
assign Simbolo[28][35] = 9'b101000000;
assign Simbolo[28][36] = 9'b100100000;
assign Simbolo[28][52] = 9'b101101001;
assign Simbolo[28][53] = 9'b100000000;
assign Simbolo[28][54] = 9'b100000000;
assign Simbolo[28][55] = 9'b100000000;
assign Simbolo[28][56] = 9'b100000000;
assign Simbolo[28][61] = 9'b100100000;
assign Simbolo[28][62] = 9'b100000000;
assign Simbolo[28][63] = 9'b100000000;
assign Simbolo[29][7] = 9'b100000000;
assign Simbolo[29][8] = 9'b100000000;
assign Simbolo[29][9] = 9'b100100000;
assign Simbolo[29][16] = 9'b100000000;
assign Simbolo[29][17] = 9'b100100100;
assign Simbolo[29][18] = 9'b101101000;
assign Simbolo[29][34] = 9'b100100000;
assign Simbolo[29][35] = 9'b101000000;
assign Simbolo[29][51] = 9'b101101001;
assign Simbolo[29][52] = 9'b100100100;
assign Simbolo[29][53] = 9'b100000000;
assign Simbolo[29][60] = 9'b101000000;
assign Simbolo[29][61] = 9'b100000000;
assign Simbolo[29][62] = 9'b100000000;
assign Simbolo[30][8] = 9'b100000000;
assign Simbolo[30][9] = 9'b100000000;
assign Simbolo[30][10] = 9'b100000000;
assign Simbolo[30][51] = 9'b101000100;
assign Simbolo[30][59] = 9'b100100000;
assign Simbolo[30][60] = 9'b100000000;
assign Simbolo[30][61] = 9'b100000000;
assign Simbolo[31][10] = 9'b100000000;
assign Simbolo[31][11] = 9'b100000000;
assign Simbolo[31][58] = 9'b100000000;
assign Simbolo[31][59] = 9'b100000000;
assign Simbolo[32][12] = 9'b100100000;
assign Simbolo[32][57] = 9'b100100000;
assign Simbolo[32][58] = 9'b100000000;
//Total de Lineas = 983

endmodule
