`timescale 1ns / 1ps

module Obs(
input enable,
input clock,
input [9:0] X, Y,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg imagen);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= X & hcount < X + RESOLUCION_X & vcount >= Y & vcount < Y + RESOLUCION_Y)
		begin
			if (Obs[vcount - Y][hcount - X][8] == 1'b1)
			begin
				red   <= Obs[vcount- Y][hcount- X][7:5];
				green <= Obs[vcount- Y][hcount- X][4:2];
            blue 	<= Obs[vcount- Y][hcount- X][1:0];
				imagen  <= 1'b1;
			end
			else
				imagen <= 0;
			end
		else
		imagen <= 0;
	end
end

parameter RESOLUCION_X = 32;
parameter RESOLUCION_Y = 15;
wire [8:0] Obs[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign Obs[0][1] = 9'b111110100;
assign Obs[0][2] = 9'b111111100;
assign Obs[0][3] = 9'b111110100;
assign Obs[0][4] = 9'b111110100;
assign Obs[0][5] = 9'b111110100;
assign Obs[0][6] = 9'b111110100;
assign Obs[0][7] = 9'b111110100;
assign Obs[0][8] = 9'b111110100;
assign Obs[0][9] = 9'b111110100;
assign Obs[0][10] = 9'b111111100;
assign Obs[0][11] = 9'b111110100;
assign Obs[0][20] = 9'b111110100;
assign Obs[0][21] = 9'b111111100;
assign Obs[0][22] = 9'b111110100;
assign Obs[0][23] = 9'b111110100;
assign Obs[0][24] = 9'b111110100;
assign Obs[0][25] = 9'b111110100;
assign Obs[0][26] = 9'b111110100;
assign Obs[0][27] = 9'b111110100;
assign Obs[0][28] = 9'b111110100;
assign Obs[0][29] = 9'b111111100;
assign Obs[0][30] = 9'b110110000;
assign Obs[1][0] = 9'b111110100;
assign Obs[1][1] = 9'b101001000;
assign Obs[1][2] = 9'b100100100;
assign Obs[1][3] = 9'b101000100;
assign Obs[1][4] = 9'b101000100;
assign Obs[1][5] = 9'b101000100;
assign Obs[1][6] = 9'b101000100;
assign Obs[1][7] = 9'b101000100;
assign Obs[1][8] = 9'b101000100;
assign Obs[1][9] = 9'b101000100;
assign Obs[1][10] = 9'b100100100;
assign Obs[1][11] = 9'b101001000;
assign Obs[1][12] = 9'b111110000;
assign Obs[1][13] = 9'b100000000;
assign Obs[1][14] = 9'b110110000;
assign Obs[1][15] = 9'b101001000;
assign Obs[1][16] = 9'b101001000;
assign Obs[1][17] = 9'b110110000;
assign Obs[1][18] = 9'b100000000;
assign Obs[1][19] = 9'b110110000;
assign Obs[1][20] = 9'b101001000;
assign Obs[1][21] = 9'b100100100;
assign Obs[1][22] = 9'b101000100;
assign Obs[1][23] = 9'b101000100;
assign Obs[1][24] = 9'b101000100;
assign Obs[1][25] = 9'b101000100;
assign Obs[1][26] = 9'b101000100;
assign Obs[1][27] = 9'b101000100;
assign Obs[1][28] = 9'b101000100;
assign Obs[1][29] = 9'b100100100;
assign Obs[1][30] = 9'b101001000;
assign Obs[1][31] = 9'b110110000;
assign Obs[2][0] = 9'b110110000;
assign Obs[2][1] = 9'b110001100;
assign Obs[2][2] = 9'b101000100;
assign Obs[2][3] = 9'b100000000;
assign Obs[2][4] = 9'b100000000;
assign Obs[2][5] = 9'b100000000;
assign Obs[2][6] = 9'b100000000;
assign Obs[2][7] = 9'b100000000;
assign Obs[2][8] = 9'b100000000;
assign Obs[2][9] = 9'b100000000;
assign Obs[2][10] = 9'b100000000;
assign Obs[2][11] = 9'b100100100;
assign Obs[2][12] = 9'b111111100;
assign Obs[2][13] = 9'b110001100;
assign Obs[2][14] = 9'b101101000;
assign Obs[2][15] = 9'b101101100;
assign Obs[2][16] = 9'b101101100;
assign Obs[2][17] = 9'b101101000;
assign Obs[2][18] = 9'b110001100;
assign Obs[2][19] = 9'b111111100;
assign Obs[2][20] = 9'b100100100;
assign Obs[2][21] = 9'b100000000;
assign Obs[2][22] = 9'b100000000;
assign Obs[2][23] = 9'b100000000;
assign Obs[2][24] = 9'b100000000;
assign Obs[2][25] = 9'b100000000;
assign Obs[2][26] = 9'b100000000;
assign Obs[2][27] = 9'b100000000;
assign Obs[2][28] = 9'b100000000;
assign Obs[2][29] = 9'b101000100;
assign Obs[2][30] = 9'b110001100;
assign Obs[2][31] = 9'b110110000;
assign Obs[3][1] = 9'b111111100;
assign Obs[3][2] = 9'b110001100;
assign Obs[3][3] = 9'b101001000;
assign Obs[3][4] = 9'b100000000;
assign Obs[3][5] = 9'b100100100;
assign Obs[3][6] = 9'b100100100;
assign Obs[3][7] = 9'b100100100;
assign Obs[3][8] = 9'b100100100;
assign Obs[3][9] = 9'b100100100;
assign Obs[3][10] = 9'b100100100;
assign Obs[3][11] = 9'b100100100;
assign Obs[3][12] = 9'b101101100;
assign Obs[3][13] = 9'b111111100;
assign Obs[3][14] = 9'b101000100;
assign Obs[3][15] = 9'b101001000;
assign Obs[3][16] = 9'b101001000;
assign Obs[3][17] = 9'b101000100;
assign Obs[3][18] = 9'b111111100;
assign Obs[3][19] = 9'b101101100;
assign Obs[3][20] = 9'b100100100;
assign Obs[3][21] = 9'b100100100;
assign Obs[3][22] = 9'b100100100;
assign Obs[3][23] = 9'b100100100;
assign Obs[3][24] = 9'b100100100;
assign Obs[3][25] = 9'b100100100;
assign Obs[3][26] = 9'b100100100;
assign Obs[3][27] = 9'b100000000;
assign Obs[3][28] = 9'b101001000;
assign Obs[3][29] = 9'b110001100;
assign Obs[3][30] = 9'b111110100;
assign Obs[4][2] = 9'b111110100;
assign Obs[4][3] = 9'b110010000;
assign Obs[4][4] = 9'b101001000;
assign Obs[4][5] = 9'b100100100;
assign Obs[4][6] = 9'b100100100;
assign Obs[4][7] = 9'b100100100;
assign Obs[4][8] = 9'b100100100;
assign Obs[4][9] = 9'b100100100;
assign Obs[4][10] = 9'b100100100;
assign Obs[4][11] = 9'b100100000;
assign Obs[4][12] = 9'b100000000;
assign Obs[4][13] = 9'b101101100;
assign Obs[4][14] = 9'b100100100;
assign Obs[4][15] = 9'b100000000;
assign Obs[4][16] = 9'b100000000;
assign Obs[4][17] = 9'b100100100;
assign Obs[4][18] = 9'b101101100;
assign Obs[4][19] = 9'b100000000;
assign Obs[4][20] = 9'b100100000;
assign Obs[4][21] = 9'b100100100;
assign Obs[4][22] = 9'b100100100;
assign Obs[4][23] = 9'b100100100;
assign Obs[4][24] = 9'b100100100;
assign Obs[4][25] = 9'b100100100;
assign Obs[4][26] = 9'b100100100;
assign Obs[4][27] = 9'b101001000;
assign Obs[4][28] = 9'b110010000;
assign Obs[4][29] = 9'b110010000;
assign Obs[5][3] = 9'b111111100;
assign Obs[5][4] = 9'b110110000;
assign Obs[5][5] = 9'b100000000;
assign Obs[5][6] = 9'b100100100;
assign Obs[5][7] = 9'b100100100;
assign Obs[5][8] = 9'b100100100;
assign Obs[5][9] = 9'b100100100;
assign Obs[5][10] = 9'b100100100;
assign Obs[5][11] = 9'b100100100;
assign Obs[5][12] = 9'b100100100;
assign Obs[5][13] = 9'b100000000;
assign Obs[5][14] = 9'b100100000;
assign Obs[5][15] = 9'b100100100;
assign Obs[5][16] = 9'b100100100;
assign Obs[5][17] = 9'b100100000;
assign Obs[5][18] = 9'b100000000;
assign Obs[5][19] = 9'b100100100;
assign Obs[5][20] = 9'b100100100;
assign Obs[5][21] = 9'b100100100;
assign Obs[5][22] = 9'b100100100;
assign Obs[5][23] = 9'b100100100;
assign Obs[5][24] = 9'b100100100;
assign Obs[5][25] = 9'b100100100;
assign Obs[5][26] = 9'b100000000;
assign Obs[5][27] = 9'b110110000;
assign Obs[5][28] = 9'b111110100;
assign Obs[6][3] = 9'b111111100;
assign Obs[6][4] = 9'b110110000;
assign Obs[6][5] = 9'b100000000;
assign Obs[6][6] = 9'b100100100;
assign Obs[6][7] = 9'b100100100;
assign Obs[6][8] = 9'b100100100;
assign Obs[6][9] = 9'b100100100;
assign Obs[6][10] = 9'b100100100;
assign Obs[6][11] = 9'b100100100;
assign Obs[6][12] = 9'b100100100;
assign Obs[6][13] = 9'b100100100;
assign Obs[6][14] = 9'b100100100;
assign Obs[6][15] = 9'b100100100;
assign Obs[6][16] = 9'b100100100;
assign Obs[6][17] = 9'b100100100;
assign Obs[6][18] = 9'b100100100;
assign Obs[6][19] = 9'b100100100;
assign Obs[6][20] = 9'b100100100;
assign Obs[6][21] = 9'b100100100;
assign Obs[6][22] = 9'b100100100;
assign Obs[6][23] = 9'b100100100;
assign Obs[6][24] = 9'b100100100;
assign Obs[6][25] = 9'b100100100;
assign Obs[6][26] = 9'b100000000;
assign Obs[6][27] = 9'b110110000;
assign Obs[6][28] = 9'b111111100;
assign Obs[7][4] = 9'b110010000;
assign Obs[7][5] = 9'b100100100;
assign Obs[7][6] = 9'b100100100;
assign Obs[7][7] = 9'b100100100;
assign Obs[7][8] = 9'b100100100;
assign Obs[7][9] = 9'b100100100;
assign Obs[7][10] = 9'b100100100;
assign Obs[7][11] = 9'b100100100;
assign Obs[7][12] = 9'b100100100;
assign Obs[7][13] = 9'b100100100;
assign Obs[7][14] = 9'b100100100;
assign Obs[7][15] = 9'b100100100;
assign Obs[7][16] = 9'b100100100;
assign Obs[7][17] = 9'b100100100;
assign Obs[7][18] = 9'b100100100;
assign Obs[7][19] = 9'b100100100;
assign Obs[7][20] = 9'b100100100;
assign Obs[7][21] = 9'b100100100;
assign Obs[7][22] = 9'b100100100;
assign Obs[7][23] = 9'b100100100;
assign Obs[7][24] = 9'b100100100;
assign Obs[7][25] = 9'b100100100;
assign Obs[7][26] = 9'b100100100;
assign Obs[7][27] = 9'b110010000;
assign Obs[7][28] = 9'b111111100;
assign Obs[8][5] = 9'b110110000;
assign Obs[8][6] = 9'b110110000;
assign Obs[8][7] = 9'b111110000;
assign Obs[8][8] = 9'b101001000;
assign Obs[8][9] = 9'b100000000;
assign Obs[8][10] = 9'b100000000;
assign Obs[8][11] = 9'b100100100;
assign Obs[8][12] = 9'b100100100;
assign Obs[8][13] = 9'b100100100;
assign Obs[8][14] = 9'b100100100;
assign Obs[8][15] = 9'b100100100;
assign Obs[8][16] = 9'b100100100;
assign Obs[8][17] = 9'b100100100;
assign Obs[8][18] = 9'b100100100;
assign Obs[8][19] = 9'b100100100;
assign Obs[8][20] = 9'b100100100;
assign Obs[8][21] = 9'b100000000;
assign Obs[8][22] = 9'b100000000;
assign Obs[8][23] = 9'b101001000;
assign Obs[8][24] = 9'b111110100;
assign Obs[8][25] = 9'b110110000;
assign Obs[8][26] = 9'b110110000;
assign Obs[8][27] = 9'b110010000;
assign Obs[9][8] = 9'b110010000;
assign Obs[9][9] = 9'b111110000;
assign Obs[9][10] = 9'b101101100;
assign Obs[9][11] = 9'b100000000;
assign Obs[9][12] = 9'b100000000;
assign Obs[9][13] = 9'b100100100;
assign Obs[9][14] = 9'b100100100;
assign Obs[9][15] = 9'b100100100;
assign Obs[9][16] = 9'b100100100;
assign Obs[9][17] = 9'b100100100;
assign Obs[9][18] = 9'b100100100;
assign Obs[9][19] = 9'b100000000;
assign Obs[9][20] = 9'b100000000;
assign Obs[9][21] = 9'b101101100;
assign Obs[9][22] = 9'b111110000;
assign Obs[9][23] = 9'b110010000;
assign Obs[10][8] = 9'b110110000;
assign Obs[10][9] = 9'b111111100;
assign Obs[10][10] = 9'b110010000;
assign Obs[10][11] = 9'b110010000;
assign Obs[10][12] = 9'b110001100;
assign Obs[10][13] = 9'b100100100;
assign Obs[10][14] = 9'b100000000;
assign Obs[10][15] = 9'b100100100;
assign Obs[10][16] = 9'b100100100;
assign Obs[10][17] = 9'b100000000;
assign Obs[10][18] = 9'b100100100;
assign Obs[10][19] = 9'b110001100;
assign Obs[10][20] = 9'b110010000;
assign Obs[10][21] = 9'b110001100;
assign Obs[10][22] = 9'b111111100;
assign Obs[11][11] = 9'b111111100;
assign Obs[11][12] = 9'b111111100;
assign Obs[11][13] = 9'b101101100;
assign Obs[11][14] = 9'b100100100;
assign Obs[11][15] = 9'b100000000;
assign Obs[11][16] = 9'b100000000;
assign Obs[11][17] = 9'b100100100;
assign Obs[11][18] = 9'b101101100;
assign Obs[11][19] = 9'b111110100;
assign Obs[11][20] = 9'b111111100;
assign Obs[12][13] = 9'b111111100;
assign Obs[12][14] = 9'b101101100;
assign Obs[12][15] = 9'b100100100;
assign Obs[12][16] = 9'b100100100;
assign Obs[12][17] = 9'b101101100;
assign Obs[12][18] = 9'b111111100;
assign Obs[13][14] = 9'b111111100;
assign Obs[13][15] = 9'b101101100;
assign Obs[13][16] = 9'b101101000;
assign Obs[13][17] = 9'b111111100;
assign Obs[14][15] = 9'b110110000;
assign Obs[14][16] = 9'b110110000;
//Total de Lineas = 297
endmodule