`timescale 1ns / 1ps

module Obs2(
input enable,
input clock,
input [9:0] X, Y,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg imagen);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= X & hcount < X + RESOLUCION_X & vcount >= Y & vcount < Y + RESOLUCION_Y)
		begin
			if (Acertijo[vcount - Y][hcount - X][8] == 1'b1)
			begin
				red   <= Acertijo[vcount- Y][hcount- X][7:5];
				green <= Acertijo[vcount- Y][hcount- X][4:2];
            blue 	<= Acertijo[vcount- Y][hcount- X][1:0];
				imagen  <= 1'b1;
			end
			else
				imagen <= 0;
			end
		else
		imagen <= 0;
	end
end

parameter RESOLUCION_X = 20;
parameter RESOLUCION_Y = 32;
wire [8:0] Acertijo[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign Acertijo[0][5] = 9'b100100100;
assign Acertijo[0][6] = 9'b100100100;
assign Acertijo[0][7] = 9'b100100100;
assign Acertijo[0][8] = 9'b100100100;
assign Acertijo[0][9] = 9'b100100100;
assign Acertijo[0][10] = 9'b100100100;
assign Acertijo[0][11] = 9'b100100100;
assign Acertijo[0][12] = 9'b100100000;
assign Acertijo[1][4] = 9'b100100000;
assign Acertijo[1][5] = 9'b100100100;
assign Acertijo[1][6] = 9'b100101100;
assign Acertijo[1][7] = 9'b100111100;
assign Acertijo[1][8] = 9'b100111100;
assign Acertijo[1][9] = 9'b100111100;
assign Acertijo[1][10] = 9'b100111100;
assign Acertijo[1][11] = 9'b100110100;
assign Acertijo[1][12] = 9'b100101000;
assign Acertijo[1][13] = 9'b100100100;
assign Acertijo[1][14] = 9'b100100000;
assign Acertijo[2][3] = 9'b100100000;
assign Acertijo[2][4] = 9'b100101000;
assign Acertijo[2][5] = 9'b100110000;
assign Acertijo[2][6] = 9'b100101100;
assign Acertijo[2][7] = 9'b100101100;
assign Acertijo[2][8] = 9'b100101100;
assign Acertijo[2][9] = 9'b100101100;
assign Acertijo[2][10] = 9'b100101100;
assign Acertijo[2][11] = 9'b100110100;
assign Acertijo[2][12] = 9'b100111100;
assign Acertijo[2][13] = 9'b100110000;
assign Acertijo[2][14] = 9'b100101000;
assign Acertijo[2][15] = 9'b100100100;
assign Acertijo[3][2] = 9'b100100000;
assign Acertijo[3][3] = 9'b100101000;
assign Acertijo[3][4] = 9'b100111100;
assign Acertijo[3][5] = 9'b100100100;
assign Acertijo[3][6] = 9'b100100000;
assign Acertijo[3][7] = 9'b100100000;
assign Acertijo[3][8] = 9'b100100000;
assign Acertijo[3][9] = 9'b100100000;
assign Acertijo[3][10] = 9'b100100000;
assign Acertijo[3][11] = 9'b100101000;
assign Acertijo[3][12] = 9'b100111100;
assign Acertijo[3][13] = 9'b100111100;
assign Acertijo[3][14] = 9'b100111100;
assign Acertijo[3][15] = 9'b100101100;
assign Acertijo[3][16] = 9'b100100100;
assign Acertijo[4][1] = 9'b100100000;
assign Acertijo[4][2] = 9'b100101000;
assign Acertijo[4][3] = 9'b100110100;
assign Acertijo[4][4] = 9'b100100100;
assign Acertijo[4][5] = 9'b100100000;
assign Acertijo[4][6] = 9'b100100100;
assign Acertijo[4][7] = 9'b100100100;
assign Acertijo[4][8] = 9'b100100100;
assign Acertijo[4][9] = 9'b100100100;
assign Acertijo[4][10] = 9'b100100100;
assign Acertijo[4][11] = 9'b100100000;
assign Acertijo[4][12] = 9'b100001000;
assign Acertijo[4][13] = 9'b100110000;
assign Acertijo[4][14] = 9'b100111100;
assign Acertijo[4][15] = 9'b100110100;
assign Acertijo[4][16] = 9'b100100100;
assign Acertijo[5][1] = 9'b100100000;
assign Acertijo[5][2] = 9'b100101100;
assign Acertijo[5][3] = 9'b100111100;
assign Acertijo[5][4] = 9'b100101100;
assign Acertijo[5][5] = 9'b100100000;
assign Acertijo[5][6] = 9'b100100100;
assign Acertijo[5][7] = 9'b100100100;
assign Acertijo[5][8] = 9'b100000100;
assign Acertijo[5][9] = 9'b100100100;
assign Acertijo[5][10] = 9'b100100100;
assign Acertijo[5][11] = 9'b100100100;
assign Acertijo[5][12] = 9'b101100101;
assign Acertijo[5][13] = 9'b101000100;
assign Acertijo[5][14] = 9'b100010000;
assign Acertijo[5][15] = 9'b100111100;
assign Acertijo[5][16] = 9'b100101100;
assign Acertijo[5][17] = 9'b100100000;
assign Acertijo[6][1] = 9'b100100000;
assign Acertijo[6][2] = 9'b100101100;
assign Acertijo[6][3] = 9'b100111100;
assign Acertijo[6][4] = 9'b100111100;
assign Acertijo[6][5] = 9'b100101000;
assign Acertijo[6][6] = 9'b100100000;
assign Acertijo[6][7] = 9'b100100100;
assign Acertijo[6][8] = 9'b110001010;
assign Acertijo[6][9] = 9'b110101011;
assign Acertijo[6][11] = 9'b110101011;
assign Acertijo[6][12] = 9'b110101011;
assign Acertijo[6][13] = 9'b110000110;
assign Acertijo[6][14] = 9'b101101001;
assign Acertijo[6][15] = 9'b110001010;
assign Acertijo[6][16] = 9'b101101101;
assign Acertijo[6][17] = 9'b100101100;
assign Acertijo[6][18] = 9'b100100000;
assign Acertijo[6][19] = 9'b100100100;
assign Acertijo[7][1] = 9'b100000000;
assign Acertijo[7][2] = 9'b100101100;
assign Acertijo[7][3] = 9'b100111100;
assign Acertijo[7][4] = 9'b100111100;
assign Acertijo[7][5] = 9'b100101100;
assign Acertijo[7][6] = 9'b100100000;
assign Acertijo[7][7] = 9'b110000101;
assign Acertijo[7][8] = 9'b110000110;
assign Acertijo[7][9] = 9'b100100100;
assign Acertijo[7][10] = 9'b100100100;
assign Acertijo[7][11] = 9'b100100100;
assign Acertijo[7][12] = 9'b110001010;
assign Acertijo[7][13] = 9'b110001011;
assign Acertijo[7][14] = 9'b110001011;
assign Acertijo[7][15] = 9'b110000111;
assign Acertijo[7][16] = 9'b110001011;
assign Acertijo[7][17] = 9'b110001010;
assign Acertijo[7][18] = 9'b110000110;
assign Acertijo[7][19] = 9'b100100100;
assign Acertijo[8][1] = 9'b100000000;
assign Acertijo[8][2] = 9'b100101100;
assign Acertijo[8][3] = 9'b100111100;
assign Acertijo[8][4] = 9'b100111100;
assign Acertijo[8][5] = 9'b100001100;
assign Acertijo[8][6] = 9'b101100101;
assign Acertijo[8][7] = 9'b110001010;
assign Acertijo[8][8] = 9'b100100100;
assign Acertijo[8][9] = 9'b100100100;
assign Acertijo[8][10] = 9'b100100100;
assign Acertijo[8][11] = 9'b100100100;
assign Acertijo[8][12] = 9'b110001010;
assign Acertijo[8][13] = 9'b110001011;
assign Acertijo[8][14] = 9'b110001011;
assign Acertijo[8][15] = 9'b110001011;
assign Acertijo[8][16] = 9'b110001010;
assign Acertijo[8][17] = 9'b110001010;
assign Acertijo[8][18] = 9'b101000101;
assign Acertijo[8][19] = 9'b100000000;
assign Acertijo[9][1] = 9'b100000000;
assign Acertijo[9][2] = 9'b100000000;
assign Acertijo[9][3] = 9'b100001100;
assign Acertijo[9][4] = 9'b100001100;
assign Acertijo[9][5] = 9'b100000000;
assign Acertijo[9][6] = 9'b101100101;
assign Acertijo[9][7] = 9'b101000100;
assign Acertijo[9][8] = 9'b100000000;
assign Acertijo[9][9] = 9'b100000100;
assign Acertijo[9][10] = 9'b100000000;
assign Acertijo[9][11] = 9'b100100100;
assign Acertijo[9][12] = 9'b110001010;
assign Acertijo[9][13] = 9'b110101011;
assign Acertijo[9][14] = 9'b110000110;
assign Acertijo[9][15] = 9'b101101001;
assign Acertijo[9][16] = 9'b100111100;
assign Acertijo[9][17] = 9'b100101100;
assign Acertijo[9][18] = 9'b100100000;
assign Acertijo[10][0] = 9'b100000000;
assign Acertijo[10][1] = 9'b100100100;
assign Acertijo[10][2] = 9'b101000100;
assign Acertijo[10][3] = 9'b101000101;
assign Acertijo[10][4] = 9'b101000101;
assign Acertijo[10][5] = 9'b101100101;
assign Acertijo[10][6] = 9'b111101011;
assign Acertijo[10][7] = 9'b101000101;
assign Acertijo[10][8] = 9'b100100100;
assign Acertijo[10][9] = 9'b101000101;
assign Acertijo[10][10] = 9'b100100100;
assign Acertijo[10][11] = 9'b110001010;
assign Acertijo[10][12] = 9'b110101011;
assign Acertijo[10][13] = 9'b110000110;
assign Acertijo[10][14] = 9'b100100100;
assign Acertijo[10][15] = 9'b100010000;
assign Acertijo[10][16] = 9'b100110100;
assign Acertijo[10][17] = 9'b100101000;
assign Acertijo[10][18] = 9'b100100000;
assign Acertijo[11][0] = 9'b100100100;
assign Acertijo[11][1] = 9'b101100101;
assign Acertijo[11][2] = 9'b110101011;
assign Acertijo[11][3] = 9'b101100101;
assign Acertijo[11][4] = 9'b101100101;
assign Acertijo[11][5] = 9'b110001010;
assign Acertijo[11][6] = 9'b101000101;
assign Acertijo[11][7] = 9'b110001011;
assign Acertijo[11][8] = 9'b110101011;
assign Acertijo[11][9] = 9'b110101011;
assign Acertijo[11][10] = 9'b110101011;
assign Acertijo[11][11] = 9'b110101011;
assign Acertijo[11][12] = 9'b101100101;
assign Acertijo[11][13] = 9'b101000101;
assign Acertijo[11][14] = 9'b100010000;
assign Acertijo[11][15] = 9'b100111100;
assign Acertijo[11][16] = 9'b100110000;
assign Acertijo[11][17] = 9'b100100000;
assign Acertijo[12][0] = 9'b100100100;
assign Acertijo[12][1] = 9'b101100101;
assign Acertijo[12][2] = 9'b110101011;
assign Acertijo[12][3] = 9'b100100100;
assign Acertijo[12][4] = 9'b100100100;
assign Acertijo[12][5] = 9'b101100101;
assign Acertijo[12][6] = 9'b100000000;
assign Acertijo[12][7] = 9'b101000101;
assign Acertijo[12][8] = 9'b101000101;
assign Acertijo[12][9] = 9'b101000101;
assign Acertijo[12][10] = 9'b101000101;
assign Acertijo[12][11] = 9'b101000101;
assign Acertijo[12][12] = 9'b100001000;
assign Acertijo[12][13] = 9'b100110000;
assign Acertijo[12][14] = 9'b100111100;
assign Acertijo[12][15] = 9'b100111100;
assign Acertijo[12][16] = 9'b100110000;
assign Acertijo[12][17] = 9'b100100000;
assign Acertijo[13][0] = 9'b100000100;
assign Acertijo[13][1] = 9'b100100100;
assign Acertijo[13][2] = 9'b110001010;
assign Acertijo[13][3] = 9'b101100101;
assign Acertijo[13][4] = 9'b101000100;
assign Acertijo[13][5] = 9'b101100101;
assign Acertijo[13][6] = 9'b100000100;
assign Acertijo[13][7] = 9'b100000100;
assign Acertijo[13][8] = 9'b100000000;
assign Acertijo[13][9] = 9'b100000000;
assign Acertijo[13][10] = 9'b100000000;
assign Acertijo[13][11] = 9'b100001100;
assign Acertijo[13][12] = 9'b100111100;
assign Acertijo[13][13] = 9'b100111100;
assign Acertijo[13][14] = 9'b100110100;
assign Acertijo[13][15] = 9'b100110100;
assign Acertijo[13][16] = 9'b100101000;
assign Acertijo[13][17] = 9'b100100000;
assign Acertijo[14][1] = 9'b100000000;
assign Acertijo[14][2] = 9'b100100100;
assign Acertijo[14][3] = 9'b110001010;
assign Acertijo[14][4] = 9'b110001010;
assign Acertijo[14][5] = 9'b101100101;
assign Acertijo[14][6] = 9'b100000100;
assign Acertijo[14][7] = 9'b100100100;
assign Acertijo[14][8] = 9'b100100000;
assign Acertijo[14][9] = 9'b100101000;
assign Acertijo[14][10] = 9'b100110000;
assign Acertijo[14][11] = 9'b100110100;
assign Acertijo[14][12] = 9'b100110100;
assign Acertijo[14][13] = 9'b100110100;
assign Acertijo[14][14] = 9'b100110100;
assign Acertijo[14][15] = 9'b100101000;
assign Acertijo[14][16] = 9'b100100000;
assign Acertijo[15][2] = 9'b100000100;
assign Acertijo[15][3] = 9'b110001010;
assign Acertijo[15][4] = 9'b110101011;
assign Acertijo[15][5] = 9'b101100101;
assign Acertijo[15][6] = 9'b100000000;
assign Acertijo[15][7] = 9'b100100100;
assign Acertijo[15][8] = 9'b100110000;
assign Acertijo[15][9] = 9'b100110100;
assign Acertijo[15][10] = 9'b100111100;
assign Acertijo[15][11] = 9'b100111100;
assign Acertijo[15][12] = 9'b100110100;
assign Acertijo[15][13] = 9'b100110100;
assign Acertijo[15][14] = 9'b100101100;
assign Acertijo[15][15] = 9'b100100000;
assign Acertijo[16][2] = 9'b100000100;
assign Acertijo[16][3] = 9'b101101001;
assign Acertijo[16][4] = 9'b101100101;
assign Acertijo[16][5] = 9'b100100100;
assign Acertijo[16][6] = 9'b100100100;
assign Acertijo[16][7] = 9'b100110000;
assign Acertijo[16][8] = 9'b100111100;
assign Acertijo[16][9] = 9'b100111100;
assign Acertijo[16][10] = 9'b100110000;
assign Acertijo[16][11] = 9'b100110000;
assign Acertijo[16][12] = 9'b100110000;
assign Acertijo[16][13] = 9'b100100100;
assign Acertijo[16][14] = 9'b100100100;
assign Acertijo[17][2] = 9'b100100100;
assign Acertijo[17][3] = 9'b100100100;
assign Acertijo[17][4] = 9'b100100000;
assign Acertijo[17][5] = 9'b100100000;
assign Acertijo[17][6] = 9'b100101100;
assign Acertijo[17][7] = 9'b100111100;
assign Acertijo[17][8] = 9'b100110100;
assign Acertijo[17][9] = 9'b100110000;
assign Acertijo[17][10] = 9'b100101000;
assign Acertijo[17][11] = 9'b100100000;
assign Acertijo[17][12] = 9'b100100100;
assign Acertijo[17][13] = 9'b100000000;
assign Acertijo[18][5] = 9'b100100100;
assign Acertijo[18][6] = 9'b100110000;
assign Acertijo[18][7] = 9'b100111100;
assign Acertijo[18][8] = 9'b100101100;
assign Acertijo[18][9] = 9'b100100000;
assign Acertijo[18][10] = 9'b100100100;
assign Acertijo[19][5] = 9'b100101000;
assign Acertijo[19][6] = 9'b100111100;
assign Acertijo[19][7] = 9'b100110100;
assign Acertijo[19][8] = 9'b100100100;
assign Acertijo[19][9] = 9'b100100000;
assign Acertijo[19][10] = 9'b100100100;
assign Acertijo[19][11] = 9'b100100000;
assign Acertijo[19][12] = 9'b100000000;
assign Acertijo[20][5] = 9'b100101000;
assign Acertijo[20][6] = 9'b100111100;
assign Acertijo[20][7] = 9'b100101100;
assign Acertijo[20][8] = 9'b100100100;
assign Acertijo[20][9] = 9'b100100100;
assign Acertijo[20][10] = 9'b100100000;
assign Acertijo[20][11] = 9'b100101000;
assign Acertijo[20][12] = 9'b100100100;
assign Acertijo[21][5] = 9'b100101000;
assign Acertijo[21][6] = 9'b100111100;
assign Acertijo[21][7] = 9'b100101100;
assign Acertijo[21][8] = 9'b100100000;
assign Acertijo[21][9] = 9'b100100000;
assign Acertijo[21][10] = 9'b100101000;
assign Acertijo[21][11] = 9'b100110100;
assign Acertijo[21][12] = 9'b100100100;
assign Acertijo[22][5] = 9'b100100100;
assign Acertijo[22][6] = 9'b100110000;
assign Acertijo[22][7] = 9'b100111100;
assign Acertijo[22][8] = 9'b100110000;
assign Acertijo[22][9] = 9'b100110000;
assign Acertijo[22][10] = 9'b100110100;
assign Acertijo[22][11] = 9'b100110100;
assign Acertijo[22][12] = 9'b100100100;
assign Acertijo[23][5] = 9'b100100000;
assign Acertijo[23][6] = 9'b100100100;
assign Acertijo[23][7] = 9'b100110000;
assign Acertijo[23][8] = 9'b100110100;
assign Acertijo[23][9] = 9'b100110100;
assign Acertijo[23][10] = 9'b100110100;
assign Acertijo[23][11] = 9'b100101000;
assign Acertijo[23][12] = 9'b100100000;
assign Acertijo[24][6] = 9'b100100000;
assign Acertijo[24][7] = 9'b100100100;
assign Acertijo[24][8] = 9'b100100100;
assign Acertijo[24][9] = 9'b100100100;
assign Acertijo[24][10] = 9'b100100100;
assign Acertijo[24][11] = 9'b100100000;
assign Acertijo[25][6] = 9'b100100000;
assign Acertijo[25][7] = 9'b100100100;
assign Acertijo[25][8] = 9'b100110100;
assign Acertijo[25][9] = 9'b100110000;
assign Acertijo[25][10] = 9'b100100000;
assign Acertijo[25][11] = 9'b100100000;
assign Acertijo[26][5] = 9'b100100000;
assign Acertijo[26][6] = 9'b100100100;
assign Acertijo[26][7] = 9'b100110000;
assign Acertijo[26][8] = 9'b100111100;
assign Acertijo[26][9] = 9'b100111100;
assign Acertijo[26][10] = 9'b100101100;
assign Acertijo[26][11] = 9'b100100100;
assign Acertijo[27][5] = 9'b100100000;
assign Acertijo[27][6] = 9'b100101100;
assign Acertijo[27][7] = 9'b100111100;
assign Acertijo[27][8] = 9'b100110100;
assign Acertijo[27][9] = 9'b100110100;
assign Acertijo[27][10] = 9'b100111100;
assign Acertijo[27][11] = 9'b100101000;
assign Acertijo[28][5] = 9'b100100000;
assign Acertijo[28][6] = 9'b100101100;
assign Acertijo[28][7] = 9'b100111100;
assign Acertijo[28][8] = 9'b100110100;
assign Acertijo[28][9] = 9'b100110100;
assign Acertijo[28][10] = 9'b100111100;
assign Acertijo[28][11] = 9'b100101000;
assign Acertijo[29][5] = 9'b100100000;
assign Acertijo[29][6] = 9'b100101000;
assign Acertijo[29][7] = 9'b100110000;
assign Acertijo[29][8] = 9'b100110100;
assign Acertijo[29][9] = 9'b100111100;
assign Acertijo[29][10] = 9'b100101100;
assign Acertijo[29][11] = 9'b100100100;
assign Acertijo[30][6] = 9'b100100000;
assign Acertijo[30][7] = 9'b100101000;
assign Acertijo[30][8] = 9'b100110100;
assign Acertijo[30][9] = 9'b100110000;
assign Acertijo[30][10] = 9'b100100100;
assign Acertijo[30][11] = 9'b100100000;
assign Acertijo[31][7] = 9'b100100000;
assign Acertijo[31][8] = 9'b100100100;
assign Acertijo[31][9] = 9'b100100100;
assign Acertijo[31][10] = 9'b100100000;
//Total de Lineas = 378

endmodule
