`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:53:05 04/30/2021 
// Design Name: 
// Module Name:    Over 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Over(
input enable,
input clock,
input [9:0] X, Y,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg imagen);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= X & hcount < X + RESOLUCION_X & vcount >= Y & vcount < Y + RESOLUCION_Y)
		begin
			if (Over[vcount - Y][hcount - X][8] == 1'b1)
			begin
				red   <= Over[vcount- Y][hcount- X][7:5];
				green <= Over[vcount- Y][hcount- X][4:2];
            blue 	<= Over[vcount- Y][hcount- X][1:0];
				imagen  <= 1'b1;
			end
			else
				imagen <= 0;
			end
		else
		imagen <= 0;
	end
end
parameter RESOLUCION_X = 70;
parameter RESOLUCION_Y = 40;
wire [8:0] Over[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign Over[1][33] = 9'b110010001;
assign Over[1][36] = 9'b110010001;
assign Over[2][32] = 9'b110111111;
assign Over[2][33] = 9'b111111111;
assign Over[2][36] = 9'b110010001;
assign Over[3][32] = 9'b110010010;
assign Over[3][33] = 9'b110110110;
assign Over[3][36] = 9'b110010010;
assign Over[4][20] = 9'b111111111;
assign Over[4][21] = 9'b110010010;
assign Over[4][32] = 9'b110010010;
assign Over[4][35] = 9'b111111111;
assign Over[4][36] = 9'b110010010;
assign Over[4][37] = 9'b110010001;
assign Over[4][47] = 9'b110110110;
assign Over[4][48] = 9'b110110110;
assign Over[4][49] = 9'b101001000;
assign Over[5][19] = 9'b111111111;
assign Over[5][20] = 9'b110010001;
assign Over[5][21] = 9'b100100100;
assign Over[5][22] = 9'b101101101;
assign Over[5][23] = 9'b110110110;
assign Over[5][32] = 9'b111111111;
assign Over[5][33] = 9'b101001001;
assign Over[5][34] = 9'b101110001;
assign Over[5][35] = 9'b110110110;
assign Over[5][36] = 9'b101001101;
assign Over[5][37] = 9'b101101101;
assign Over[5][46] = 9'b111111111;
assign Over[5][47] = 9'b111111111;
assign Over[5][48] = 9'b101001000;
assign Over[5][49] = 9'b101001001;
assign Over[5][50] = 9'b101001001;
assign Over[6][19] = 9'b110010010;
assign Over[6][20] = 9'b100000000;
assign Over[6][21] = 9'b100000000;
assign Over[6][22] = 9'b100000100;
assign Over[6][23] = 9'b101101101;
assign Over[6][24] = 9'b111111111;
assign Over[6][32] = 9'b110110110;
assign Over[6][33] = 9'b100100100;
assign Over[6][34] = 9'b100101000;
assign Over[6][35] = 9'b100101000;
assign Over[6][36] = 9'b100100100;
assign Over[6][37] = 9'b101001001;
assign Over[6][44] = 9'b111111111;
assign Over[6][45] = 9'b111111111;
assign Over[6][46] = 9'b110010010;
assign Over[6][47] = 9'b100100100;
assign Over[6][48] = 9'b100000000;
assign Over[6][49] = 9'b100000000;
assign Over[6][50] = 9'b101110001;
assign Over[6][51] = 9'b101001001;
assign Over[7][18] = 9'b101110001;
assign Over[7][19] = 9'b100100100;
assign Over[7][20] = 9'b100000000;
assign Over[7][21] = 9'b100000000;
assign Over[7][22] = 9'b100000000;
assign Over[7][23] = 9'b100000000;
assign Over[7][24] = 9'b100100100;
assign Over[7][25] = 9'b110010001;
assign Over[7][26] = 9'b111111111;
assign Over[7][27] = 9'b111111111;
assign Over[7][32] = 9'b110010010;
assign Over[7][33] = 9'b100100100;
assign Over[7][34] = 9'b100000000;
assign Over[7][35] = 9'b100000000;
assign Over[7][36] = 9'b100000100;
assign Over[7][37] = 9'b100100100;
assign Over[7][42] = 9'b110010010;
assign Over[7][43] = 9'b110110110;
assign Over[7][44] = 9'b110010110;
assign Over[7][45] = 9'b101001001;
assign Over[7][46] = 9'b100000000;
assign Over[7][47] = 9'b100000000;
assign Over[7][48] = 9'b100000000;
assign Over[7][49] = 9'b100000000;
assign Over[7][50] = 9'b100100100;
assign Over[7][51] = 9'b110010001;
assign Over[7][52] = 9'b100100100;
assign Over[8][17] = 9'b110010010;
assign Over[8][18] = 9'b100100100;
assign Over[8][19] = 9'b100000000;
assign Over[8][20] = 9'b100000000;
assign Over[8][21] = 9'b100000000;
assign Over[8][22] = 9'b100000000;
assign Over[8][23] = 9'b100000000;
assign Over[8][24] = 9'b100000000;
assign Over[8][25] = 9'b100000000;
assign Over[8][26] = 9'b101001000;
assign Over[8][27] = 9'b110010001;
assign Over[8][28] = 9'b111111111;
assign Over[8][29] = 9'b111111111;
assign Over[8][30] = 9'b111111111;
assign Over[8][32] = 9'b110010001;
assign Over[8][33] = 9'b100000000;
assign Over[8][34] = 9'b100000000;
assign Over[8][35] = 9'b100000000;
assign Over[8][36] = 9'b100000000;
assign Over[8][37] = 9'b100100100;
assign Over[8][38] = 9'b101001001;
assign Over[8][39] = 9'b101001101;
assign Over[8][40] = 9'b101101101;
assign Over[8][41] = 9'b101110001;
assign Over[8][42] = 9'b101101101;
assign Over[8][43] = 9'b101001001;
assign Over[8][44] = 9'b100000000;
assign Over[8][45] = 9'b100000000;
assign Over[8][46] = 9'b100000000;
assign Over[8][47] = 9'b100000000;
assign Over[8][48] = 9'b100000000;
assign Over[8][49] = 9'b100000000;
assign Over[8][50] = 9'b100000000;
assign Over[8][51] = 9'b100100100;
assign Over[8][52] = 9'b101001001;
assign Over[9][16] = 9'b110111111;
assign Over[9][17] = 9'b101001001;
assign Over[9][18] = 9'b100000000;
assign Over[9][19] = 9'b100000000;
assign Over[9][20] = 9'b100000000;
assign Over[9][21] = 9'b100000000;
assign Over[9][22] = 9'b100000000;
assign Over[9][23] = 9'b100000000;
assign Over[9][24] = 9'b100000000;
assign Over[9][25] = 9'b100000000;
assign Over[9][26] = 9'b100000000;
assign Over[9][27] = 9'b100000000;
assign Over[9][28] = 9'b100100100;
assign Over[9][29] = 9'b101001001;
assign Over[9][30] = 9'b110010001;
assign Over[9][31] = 9'b110110110;
assign Over[9][32] = 9'b101101101;
assign Over[9][33] = 9'b100000000;
assign Over[9][34] = 9'b100000000;
assign Over[9][35] = 9'b100000000;
assign Over[9][36] = 9'b100000000;
assign Over[9][37] = 9'b100100100;
assign Over[9][38] = 9'b100100100;
assign Over[9][39] = 9'b100100100;
assign Over[9][40] = 9'b100100100;
assign Over[9][41] = 9'b100000000;
assign Over[9][42] = 9'b100000000;
assign Over[9][43] = 9'b100000000;
assign Over[9][44] = 9'b100000000;
assign Over[9][45] = 9'b100000000;
assign Over[9][46] = 9'b100000000;
assign Over[9][47] = 9'b100000000;
assign Over[9][48] = 9'b100000000;
assign Over[9][49] = 9'b100000000;
assign Over[9][50] = 9'b100000000;
assign Over[9][51] = 9'b100000000;
assign Over[9][52] = 9'b100100100;
assign Over[9][53] = 9'b101001000;
assign Over[10][15] = 9'b111111111;
assign Over[10][16] = 9'b101101101;
assign Over[10][17] = 9'b100000000;
assign Over[10][18] = 9'b100000000;
assign Over[10][19] = 9'b100000000;
assign Over[10][20] = 9'b100000000;
assign Over[10][21] = 9'b100000000;
assign Over[10][22] = 9'b100000000;
assign Over[10][23] = 9'b100000000;
assign Over[10][24] = 9'b100000000;
assign Over[10][25] = 9'b100000000;
assign Over[10][26] = 9'b100000000;
assign Over[10][27] = 9'b100000000;
assign Over[10][28] = 9'b100000000;
assign Over[10][29] = 9'b100000000;
assign Over[10][30] = 9'b100000000;
assign Over[10][31] = 9'b100000000;
assign Over[10][32] = 9'b100000000;
assign Over[10][33] = 9'b100000000;
assign Over[10][34] = 9'b100000000;
assign Over[10][35] = 9'b100000000;
assign Over[10][36] = 9'b100000000;
assign Over[10][37] = 9'b100000000;
assign Over[10][38] = 9'b100000000;
assign Over[10][39] = 9'b100000000;
assign Over[10][40] = 9'b100000000;
assign Over[10][41] = 9'b100000000;
assign Over[10][42] = 9'b100000000;
assign Over[10][43] = 9'b100000000;
assign Over[10][44] = 9'b100000000;
assign Over[10][45] = 9'b100000000;
assign Over[10][46] = 9'b100000000;
assign Over[10][47] = 9'b100000000;
assign Over[10][48] = 9'b100000000;
assign Over[10][49] = 9'b100000000;
assign Over[10][50] = 9'b100000000;
assign Over[10][51] = 9'b100000000;
assign Over[10][52] = 9'b100000000;
assign Over[10][53] = 9'b100101000;
assign Over[10][54] = 9'b100100100;
assign Over[11][15] = 9'b110010001;
assign Over[11][16] = 9'b100000000;
assign Over[11][17] = 9'b100000000;
assign Over[11][18] = 9'b100000000;
assign Over[11][19] = 9'b100000000;
assign Over[11][20] = 9'b100000000;
assign Over[11][21] = 9'b100000000;
assign Over[11][22] = 9'b100000000;
assign Over[11][23] = 9'b100000000;
assign Over[11][24] = 9'b100000000;
assign Over[11][25] = 9'b100000000;
assign Over[11][26] = 9'b100000000;
assign Over[11][27] = 9'b100000000;
assign Over[11][28] = 9'b100000000;
assign Over[11][29] = 9'b100000000;
assign Over[11][30] = 9'b100000000;
assign Over[11][31] = 9'b100000000;
assign Over[11][32] = 9'b100000000;
assign Over[11][33] = 9'b100000000;
assign Over[11][34] = 9'b100000000;
assign Over[11][35] = 9'b100000000;
assign Over[11][36] = 9'b100000000;
assign Over[11][37] = 9'b100000000;
assign Over[11][38] = 9'b100000000;
assign Over[11][39] = 9'b100000000;
assign Over[11][40] = 9'b100000000;
assign Over[11][41] = 9'b100000000;
assign Over[11][42] = 9'b100000000;
assign Over[11][43] = 9'b100000000;
assign Over[11][44] = 9'b100000000;
assign Over[11][45] = 9'b100000000;
assign Over[11][46] = 9'b100000000;
assign Over[11][47] = 9'b100000000;
assign Over[11][48] = 9'b100000000;
assign Over[11][49] = 9'b100000000;
assign Over[11][50] = 9'b100000000;
assign Over[11][51] = 9'b100000000;
assign Over[11][52] = 9'b100000000;
assign Over[11][53] = 9'b100000000;
assign Over[11][54] = 9'b100101000;
assign Over[11][55] = 9'b100100100;
assign Over[12][14] = 9'b110010110;
assign Over[12][15] = 9'b100100100;
assign Over[12][16] = 9'b100000000;
assign Over[12][17] = 9'b100000000;
assign Over[12][18] = 9'b100000000;
assign Over[12][19] = 9'b100000000;
assign Over[12][20] = 9'b100000000;
assign Over[12][21] = 9'b100000000;
assign Over[12][22] = 9'b100000000;
assign Over[12][23] = 9'b100000000;
assign Over[12][24] = 9'b100000000;
assign Over[12][25] = 9'b100000000;
assign Over[12][26] = 9'b100000000;
assign Over[12][27] = 9'b100000000;
assign Over[12][28] = 9'b100000000;
assign Over[12][29] = 9'b100000000;
assign Over[12][30] = 9'b100000000;
assign Over[12][31] = 9'b100000000;
assign Over[12][32] = 9'b100000000;
assign Over[12][33] = 9'b100000000;
assign Over[12][34] = 9'b100000000;
assign Over[12][35] = 9'b100000000;
assign Over[12][36] = 9'b100000000;
assign Over[12][37] = 9'b100000000;
assign Over[12][38] = 9'b100000000;
assign Over[12][39] = 9'b100000000;
assign Over[12][40] = 9'b100000000;
assign Over[12][41] = 9'b100000000;
assign Over[12][42] = 9'b100000000;
assign Over[12][43] = 9'b100000000;
assign Over[12][44] = 9'b100000000;
assign Over[12][45] = 9'b100000000;
assign Over[12][46] = 9'b100000000;
assign Over[12][47] = 9'b100000000;
assign Over[12][48] = 9'b100000000;
assign Over[12][49] = 9'b100000000;
assign Over[12][50] = 9'b100000000;
assign Over[12][51] = 9'b100000000;
assign Over[12][52] = 9'b100000000;
assign Over[12][53] = 9'b100000000;
assign Over[12][54] = 9'b100000000;
assign Over[12][55] = 9'b100100100;
assign Over[13][13] = 9'b111111111;
assign Over[13][14] = 9'b101001001;
assign Over[13][15] = 9'b100000000;
assign Over[13][16] = 9'b100000000;
assign Over[13][17] = 9'b100000000;
assign Over[13][18] = 9'b100000000;
assign Over[13][19] = 9'b100000000;
assign Over[13][20] = 9'b100000000;
assign Over[13][21] = 9'b100000000;
assign Over[13][22] = 9'b100000000;
assign Over[13][23] = 9'b100000000;
assign Over[13][24] = 9'b100000000;
assign Over[13][25] = 9'b100000000;
assign Over[13][26] = 9'b100000000;
assign Over[13][27] = 9'b100000000;
assign Over[13][28] = 9'b100000000;
assign Over[13][29] = 9'b100000000;
assign Over[13][30] = 9'b100000000;
assign Over[13][31] = 9'b100000000;
assign Over[13][32] = 9'b100000000;
assign Over[13][33] = 9'b100000000;
assign Over[13][34] = 9'b100000000;
assign Over[13][35] = 9'b100000000;
assign Over[13][36] = 9'b100000000;
assign Over[13][37] = 9'b100000000;
assign Over[13][38] = 9'b100000000;
assign Over[13][39] = 9'b100000000;
assign Over[13][40] = 9'b100000000;
assign Over[13][41] = 9'b100000000;
assign Over[13][42] = 9'b100000000;
assign Over[13][43] = 9'b100000000;
assign Over[13][44] = 9'b100000000;
assign Over[13][45] = 9'b100000000;
assign Over[13][46] = 9'b100000000;
assign Over[13][47] = 9'b100000000;
assign Over[13][48] = 9'b100000000;
assign Over[13][49] = 9'b100000000;
assign Over[13][50] = 9'b100000000;
assign Over[13][51] = 9'b100000000;
assign Over[13][52] = 9'b100000000;
assign Over[13][53] = 9'b100000000;
assign Over[13][54] = 9'b100000000;
assign Over[13][55] = 9'b100100100;
assign Over[13][56] = 9'b100100100;
assign Over[14][12] = 9'b111111111;
assign Over[14][13] = 9'b101101101;
assign Over[14][14] = 9'b100000000;
assign Over[14][15] = 9'b100100100;
assign Over[14][16] = 9'b100100100;
assign Over[14][17] = 9'b101001000;
assign Over[14][18] = 9'b100100100;
assign Over[14][19] = 9'b100100100;
assign Over[14][20] = 9'b100000000;
assign Over[14][21] = 9'b100000000;
assign Over[14][22] = 9'b100000000;
assign Over[14][23] = 9'b100000000;
assign Over[14][24] = 9'b100000000;
assign Over[14][25] = 9'b100000000;
assign Over[14][26] = 9'b100000000;
assign Over[14][27] = 9'b100000000;
assign Over[14][28] = 9'b100000000;
assign Over[14][29] = 9'b100000000;
assign Over[14][30] = 9'b100000000;
assign Over[14][31] = 9'b100000000;
assign Over[14][32] = 9'b100000000;
assign Over[14][33] = 9'b100000000;
assign Over[14][34] = 9'b100000000;
assign Over[14][35] = 9'b100000000;
assign Over[14][36] = 9'b100000000;
assign Over[14][37] = 9'b100000000;
assign Over[14][38] = 9'b100000000;
assign Over[14][39] = 9'b100000000;
assign Over[14][40] = 9'b100000000;
assign Over[14][41] = 9'b100000000;
assign Over[14][42] = 9'b100000000;
assign Over[14][43] = 9'b100000000;
assign Over[14][44] = 9'b100000000;
assign Over[14][45] = 9'b100000000;
assign Over[14][46] = 9'b100000000;
assign Over[14][47] = 9'b100000000;
assign Over[14][48] = 9'b100000000;
assign Over[14][49] = 9'b100000000;
assign Over[14][50] = 9'b101001001;
assign Over[14][51] = 9'b101001001;
assign Over[14][52] = 9'b100100100;
assign Over[14][53] = 9'b100100100;
assign Over[14][54] = 9'b100000000;
assign Over[14][55] = 9'b100000000;
assign Over[14][56] = 9'b100100100;
assign Over[14][57] = 9'b100100100;
assign Over[15][12] = 9'b110010001;
assign Over[15][13] = 9'b101101101;
assign Over[15][14] = 9'b110010001;
assign Over[15][15] = 9'b110010001;
assign Over[15][16] = 9'b101101101;
assign Over[15][17] = 9'b101101101;
assign Over[15][18] = 9'b100100100;
assign Over[15][19] = 9'b100100100;
assign Over[15][20] = 9'b100101000;
assign Over[15][21] = 9'b100000000;
assign Over[15][22] = 9'b100000000;
assign Over[15][23] = 9'b100000000;
assign Over[15][24] = 9'b100000000;
assign Over[15][25] = 9'b100000000;
assign Over[15][26] = 9'b100000000;
assign Over[15][27] = 9'b100000000;
assign Over[15][28] = 9'b100000000;
assign Over[15][29] = 9'b100000000;
assign Over[15][30] = 9'b100000000;
assign Over[15][31] = 9'b100000000;
assign Over[15][32] = 9'b100000000;
assign Over[15][33] = 9'b100000000;
assign Over[15][34] = 9'b100000000;
assign Over[15][35] = 9'b100000000;
assign Over[15][36] = 9'b100000000;
assign Over[15][37] = 9'b100000000;
assign Over[15][38] = 9'b100000000;
assign Over[15][39] = 9'b100000000;
assign Over[15][40] = 9'b100000000;
assign Over[15][41] = 9'b100000000;
assign Over[15][42] = 9'b100000000;
assign Over[15][43] = 9'b100000000;
assign Over[15][44] = 9'b100000000;
assign Over[15][45] = 9'b100000000;
assign Over[15][46] = 9'b100000000;
assign Over[15][47] = 9'b100000000;
assign Over[15][48] = 9'b100000100;
assign Over[15][49] = 9'b101101101;
assign Over[15][50] = 9'b101101101;
assign Over[15][51] = 9'b101101101;
assign Over[15][52] = 9'b101101101;
assign Over[15][53] = 9'b101101101;
assign Over[15][54] = 9'b101101101;
assign Over[15][55] = 9'b101001001;
assign Over[15][56] = 9'b100100100;
assign Over[15][57] = 9'b100100100;
assign Over[15][58] = 9'b100100100;
assign Over[16][11] = 9'b110110110;
assign Over[16][12] = 9'b110010001;
assign Over[16][13] = 9'b110010001;
assign Over[16][14] = 9'b101001001;
assign Over[16][15] = 9'b100100100;
assign Over[16][16] = 9'b100100100;
assign Over[16][17] = 9'b100000000;
assign Over[16][18] = 9'b100100100;
assign Over[16][19] = 9'b100100100;
assign Over[16][20] = 9'b100101000;
assign Over[16][21] = 9'b100100100;
assign Over[16][22] = 9'b100000000;
assign Over[16][23] = 9'b100000000;
assign Over[16][24] = 9'b100000000;
assign Over[16][25] = 9'b100000000;
assign Over[16][26] = 9'b100000000;
assign Over[16][27] = 9'b100000000;
assign Over[16][28] = 9'b100000000;
assign Over[16][29] = 9'b100000000;
assign Over[16][30] = 9'b100000000;
assign Over[16][31] = 9'b100000000;
assign Over[16][32] = 9'b100000000;
assign Over[16][33] = 9'b100000000;
assign Over[16][34] = 9'b100000000;
assign Over[16][35] = 9'b100000000;
assign Over[16][36] = 9'b100000000;
assign Over[16][37] = 9'b100000000;
assign Over[16][38] = 9'b100000000;
assign Over[16][39] = 9'b100000000;
assign Over[16][40] = 9'b100000000;
assign Over[16][41] = 9'b100000000;
assign Over[16][42] = 9'b100000000;
assign Over[16][43] = 9'b100000000;
assign Over[16][44] = 9'b100000000;
assign Over[16][45] = 9'b100000000;
assign Over[16][46] = 9'b100000000;
assign Over[16][47] = 9'b100000000;
assign Over[16][48] = 9'b101110001;
assign Over[16][49] = 9'b101001001;
assign Over[16][50] = 9'b100000000;
assign Over[16][51] = 9'b100000000;
assign Over[16][52] = 9'b100100100;
assign Over[16][53] = 9'b100100100;
assign Over[16][54] = 9'b100101000;
assign Over[16][55] = 9'b101001001;
assign Over[16][56] = 9'b101001001;
assign Over[16][57] = 9'b101101101;
assign Over[16][58] = 9'b101101101;
assign Over[17][10] = 9'b101101101;
assign Over[17][11] = 9'b101001000;
assign Over[17][12] = 9'b100000000;
assign Over[17][13] = 9'b100000000;
assign Over[17][14] = 9'b100000000;
assign Over[17][15] = 9'b100000000;
assign Over[17][16] = 9'b100000000;
assign Over[17][17] = 9'b100000000;
assign Over[17][18] = 9'b100000000;
assign Over[17][19] = 9'b100000100;
assign Over[17][20] = 9'b100100100;
assign Over[17][21] = 9'b101001000;
assign Over[17][22] = 9'b100000000;
assign Over[17][23] = 9'b100000000;
assign Over[17][24] = 9'b100000000;
assign Over[17][25] = 9'b100000000;
assign Over[17][26] = 9'b100000000;
assign Over[17][27] = 9'b100000000;
assign Over[17][28] = 9'b100000000;
assign Over[17][29] = 9'b100000000;
assign Over[17][30] = 9'b100000000;
assign Over[17][31] = 9'b100000000;
assign Over[17][32] = 9'b100000000;
assign Over[17][33] = 9'b100000000;
assign Over[17][34] = 9'b100000000;
assign Over[17][35] = 9'b100000000;
assign Over[17][36] = 9'b100000000;
assign Over[17][37] = 9'b100000000;
assign Over[17][38] = 9'b100000000;
assign Over[17][39] = 9'b100000000;
assign Over[17][40] = 9'b100000000;
assign Over[17][41] = 9'b100000000;
assign Over[17][42] = 9'b100000000;
assign Over[17][43] = 9'b100000000;
assign Over[17][44] = 9'b100000000;
assign Over[17][45] = 9'b100000000;
assign Over[17][46] = 9'b100000000;
assign Over[17][47] = 9'b100100100;
assign Over[17][48] = 9'b110010001;
assign Over[17][49] = 9'b100000000;
assign Over[17][50] = 9'b100100100;
assign Over[17][51] = 9'b100000000;
assign Over[17][52] = 9'b100000000;
assign Over[17][53] = 9'b100000000;
assign Over[17][54] = 9'b100000000;
assign Over[17][55] = 9'b100000000;
assign Over[17][56] = 9'b100000000;
assign Over[17][57] = 9'b100100100;
assign Over[17][58] = 9'b101001000;
assign Over[18][11] = 9'b100000000;
assign Over[18][12] = 9'b100000000;
assign Over[18][13] = 9'b100000000;
assign Over[18][14] = 9'b100000000;
assign Over[18][15] = 9'b100000000;
assign Over[18][16] = 9'b100000000;
assign Over[18][17] = 9'b100000000;
assign Over[18][18] = 9'b100000000;
assign Over[18][19] = 9'b100000000;
assign Over[18][20] = 9'b100000000;
assign Over[18][21] = 9'b100100100;
assign Over[18][22] = 9'b100100100;
assign Over[18][23] = 9'b100000000;
assign Over[18][24] = 9'b100000000;
assign Over[18][25] = 9'b100100100;
assign Over[18][26] = 9'b101001101;
assign Over[18][27] = 9'b101110001;
assign Over[18][28] = 9'b101001001;
assign Over[18][29] = 9'b100100100;
assign Over[18][30] = 9'b100000000;
assign Over[18][31] = 9'b100000000;
assign Over[18][32] = 9'b100000000;
assign Over[18][33] = 9'b100000000;
assign Over[18][34] = 9'b100000000;
assign Over[18][35] = 9'b100000000;
assign Over[18][36] = 9'b100000000;
assign Over[18][37] = 9'b100000000;
assign Over[18][38] = 9'b100000000;
assign Over[18][39] = 9'b100000000;
assign Over[18][40] = 9'b100100100;
assign Over[18][41] = 9'b100100100;
assign Over[18][42] = 9'b100100100;
assign Over[18][43] = 9'b100000100;
assign Over[18][44] = 9'b100000000;
assign Over[18][45] = 9'b100000000;
assign Over[18][46] = 9'b100000000;
assign Over[18][47] = 9'b101101101;
assign Over[18][48] = 9'b101001000;
assign Over[18][49] = 9'b100000000;
assign Over[18][50] = 9'b100000000;
assign Over[18][51] = 9'b100000000;
assign Over[18][53] = 9'b100000000;
assign Over[18][54] = 9'b100000000;
assign Over[18][55] = 9'b100000000;
assign Over[18][56] = 9'b100000000;
assign Over[18][57] = 9'b100000000;
assign Over[18][58] = 9'b100000000;
assign Over[19][12] = 9'b100000000;
assign Over[19][13] = 9'b100000000;
assign Over[19][14] = 9'b100000000;
assign Over[19][15] = 9'b100000000;
assign Over[19][20] = 9'b100000000;
assign Over[19][21] = 9'b100100100;
assign Over[19][22] = 9'b101001000;
assign Over[19][23] = 9'b100100100;
assign Over[19][24] = 9'b110010001;
assign Over[19][25] = 9'b110110110;
assign Over[19][26] = 9'b110010001;
assign Over[19][27] = 9'b101001101;
assign Over[19][28] = 9'b100100100;
assign Over[19][29] = 9'b100100100;
assign Over[19][30] = 9'b101001000;
assign Over[19][31] = 9'b100000000;
assign Over[19][32] = 9'b100000000;
assign Over[19][33] = 9'b100000000;
assign Over[19][34] = 9'b100000000;
assign Over[19][35] = 9'b100000000;
assign Over[19][36] = 9'b100000000;
assign Over[19][37] = 9'b100000000;
assign Over[19][38] = 9'b100100100;
assign Over[19][39] = 9'b101101101;
assign Over[19][40] = 9'b101001000;
assign Over[19][41] = 9'b100100100;
assign Over[19][42] = 9'b100100100;
assign Over[19][43] = 9'b101001001;
assign Over[19][44] = 9'b101001000;
assign Over[19][45] = 9'b100100100;
assign Over[19][46] = 9'b100100100;
assign Over[19][47] = 9'b110010001;
assign Over[19][48] = 9'b100000000;
assign Over[19][49] = 9'b100000000;
assign Over[19][55] = 9'b100000000;
assign Over[19][56] = 9'b100000000;
assign Over[19][57] = 9'b100000000;
assign Over[20][22] = 9'b101001000;
assign Over[20][23] = 9'b110110110;
assign Over[20][24] = 9'b110110110;
assign Over[20][25] = 9'b101101101;
assign Over[20][30] = 9'b100101000;
assign Over[20][31] = 9'b100101000;
assign Over[20][32] = 9'b100000000;
assign Over[20][33] = 9'b100000000;
assign Over[20][34] = 9'b100000000;
assign Over[20][35] = 9'b100000000;
assign Over[20][36] = 9'b100000000;
assign Over[20][37] = 9'b100000000;
assign Over[20][38] = 9'b110010001;
assign Over[20][39] = 9'b101001001;
assign Over[20][40] = 9'b100100100;
assign Over[20][41] = 9'b100100100;
assign Over[20][42] = 9'b100000000;
assign Over[20][44] = 9'b101001000;
assign Over[20][45] = 9'b101001001;
assign Over[20][46] = 9'b101110001;
assign Over[20][47] = 9'b101001001;
assign Over[21][31] = 9'b101001001;
assign Over[21][32] = 9'b100100100;
assign Over[21][33] = 9'b100000000;
assign Over[21][34] = 9'b100000000;
assign Over[21][35] = 9'b100000000;
assign Over[21][36] = 9'b100000000;
assign Over[21][37] = 9'b101110001;
assign Over[21][38] = 9'b101101101;
assign Over[22][32] = 9'b101001001;
assign Over[22][33] = 9'b100100100;
assign Over[22][34] = 9'b100000000;
assign Over[22][35] = 9'b100000000;
assign Over[22][36] = 9'b101001001;
assign Over[22][37] = 9'b111111111;
assign Over[23][32] = 9'b101001000;
assign Over[23][33] = 9'b101001001;
assign Over[23][34] = 9'b100000000;
assign Over[23][35] = 9'b100100100;
assign Over[23][36] = 9'b110110110;
assign Over[24][32] = 9'b100100100;
assign Over[24][33] = 9'b101001001;
assign Over[24][34] = 9'b100100100;
assign Over[24][35] = 9'b101101101;
assign Over[24][36] = 9'b111110110;
assign Over[24][48] = 9'b100100100;
assign Over[24][49] = 9'b100100100;
assign Over[24][50] = 9'b100100100;
assign Over[25][18] = 9'b101001001;
assign Over[25][19] = 9'b101101101;
assign Over[25][20] = 9'b101000100;
assign Over[25][21] = 9'b101001000;
assign Over[25][22] = 9'b110010001;
assign Over[25][23] = 9'b101101101;
assign Over[25][30] = 9'b101101101;
assign Over[25][31] = 9'b110001101;
assign Over[25][32] = 9'b101101101;
assign Over[25][33] = 9'b100100100;
assign Over[25][34] = 9'b101101101;
assign Over[25][35] = 9'b110110110;
assign Over[25][37] = 9'b100100100;
assign Over[25][38] = 9'b101101101;
assign Over[25][39] = 9'b110010001;
assign Over[25][40] = 9'b110010001;
assign Over[25][41] = 9'b101101101;
assign Over[25][44] = 9'b101001001;
assign Over[25][45] = 9'b100100100;
assign Over[25][46] = 9'b100100100;
assign Over[25][47] = 9'b101001001;
assign Over[25][48] = 9'b101001001;
assign Over[25][49] = 9'b101101101;
assign Over[25][50] = 9'b101101001;
assign Over[25][51] = 9'b101101101;
assign Over[25][52] = 9'b110001101;
assign Over[25][53] = 9'b101001000;
assign Over[26][17] = 9'b101001001;
assign Over[26][18] = 9'b110010001;
assign Over[26][19] = 9'b101101101;
assign Over[26][20] = 9'b101001000;
assign Over[26][21] = 9'b101101101;
assign Over[26][22] = 9'b110010001;
assign Over[26][23] = 9'b110001101;
assign Over[26][25] = 9'b101101101;
assign Over[26][26] = 9'b101101101;
assign Over[26][27] = 9'b101001001;
assign Over[26][28] = 9'b101101101;
assign Over[26][30] = 9'b101101101;
assign Over[26][31] = 9'b110010001;
assign Over[26][32] = 9'b101001001;
assign Over[26][33] = 9'b100000000;
assign Over[26][34] = 9'b110010001;
assign Over[26][35] = 9'b110010010;
assign Over[26][36] = 9'b100100100;
assign Over[26][37] = 9'b101101101;
assign Over[26][38] = 9'b101101101;
assign Over[26][39] = 9'b101001001;
assign Over[26][40] = 9'b101001001;
assign Over[26][41] = 9'b110010001;
assign Over[26][42] = 9'b101101101;
assign Over[26][43] = 9'b101001000;
assign Over[26][44] = 9'b101101101;
assign Over[26][45] = 9'b100100100;
assign Over[26][46] = 9'b101001000;
assign Over[26][47] = 9'b110001101;
assign Over[26][48] = 9'b110001101;
assign Over[26][49] = 9'b110010001;
assign Over[26][50] = 9'b101101101;
assign Over[26][51] = 9'b110010001;
assign Over[26][52] = 9'b110010001;
assign Over[26][53] = 9'b110010001;
assign Over[26][54] = 9'b101000100;
assign Over[27][16] = 9'b101001000;
assign Over[27][17] = 9'b110010001;
assign Over[27][18] = 9'b101001001;
assign Over[27][19] = 9'b100100100;
assign Over[27][20] = 9'b101001001;
assign Over[27][21] = 9'b110010001;
assign Over[27][22] = 9'b101101101;
assign Over[27][23] = 9'b110010001;
assign Over[27][24] = 9'b101001000;
assign Over[27][25] = 9'b101101101;
assign Over[27][26] = 9'b110010001;
assign Over[27][27] = 9'b110001101;
assign Over[27][28] = 9'b110010001;
assign Over[27][29] = 9'b100100100;
assign Over[27][30] = 9'b101101101;
assign Over[27][31] = 9'b101101101;
assign Over[27][32] = 9'b100100100;
assign Over[27][36] = 9'b101101101;
assign Over[27][37] = 9'b101101101;
assign Over[27][38] = 9'b100100100;
assign Over[27][39] = 9'b100000000;
assign Over[27][40] = 9'b100000000;
assign Over[27][41] = 9'b100100100;
assign Over[27][42] = 9'b110010001;
assign Over[27][43] = 9'b101101101;
assign Over[27][44] = 9'b101101101;
assign Over[27][45] = 9'b101001000;
assign Over[27][46] = 9'b101001001;
assign Over[27][47] = 9'b110001101;
assign Over[27][48] = 9'b110001101;
assign Over[27][49] = 9'b101101101;
assign Over[27][50] = 9'b101001000;
assign Over[27][51] = 9'b110001101;
assign Over[27][52] = 9'b101001000;
assign Over[27][53] = 9'b101101101;
assign Over[27][54] = 9'b101101101;
assign Over[28][16] = 9'b101101101;
assign Over[28][17] = 9'b101101101;
assign Over[28][18] = 9'b100100100;
assign Over[28][19] = 9'b101101001;
assign Over[28][20] = 9'b110001101;
assign Over[28][21] = 9'b110010010;
assign Over[28][22] = 9'b110010001;
assign Over[28][23] = 9'b110010001;
assign Over[28][24] = 9'b101001001;
assign Over[28][25] = 9'b101101101;
assign Over[28][26] = 9'b110010010;
assign Over[28][27] = 9'b110010010;
assign Over[28][28] = 9'b110010001;
assign Over[28][29] = 9'b101001001;
assign Over[28][30] = 9'b110010001;
assign Over[28][31] = 9'b110010010;
assign Over[28][32] = 9'b101101101;
assign Over[28][36] = 9'b110001101;
assign Over[28][37] = 9'b100100100;
assign Over[28][38] = 9'b100000000;
assign Over[28][39] = 9'b100000000;
assign Over[28][40] = 9'b100000000;
assign Over[28][41] = 9'b100000000;
assign Over[28][42] = 9'b101001000;
assign Over[28][43] = 9'b110010001;
assign Over[28][44] = 9'b110010001;
assign Over[28][45] = 9'b101101001;
assign Over[28][46] = 9'b101101101;
assign Over[28][47] = 9'b110001101;
assign Over[28][48] = 9'b110010001;
assign Over[28][49] = 9'b110010010;
assign Over[28][50] = 9'b110001101;
assign Over[28][51] = 9'b110010001;
assign Over[28][52] = 9'b101001000;
assign Over[28][53] = 9'b100100100;
assign Over[28][54] = 9'b110001101;
assign Over[28][55] = 9'b101001001;
assign Over[29][15] = 9'b100100100;
assign Over[29][16] = 9'b110001101;
assign Over[29][17] = 9'b100100100;
assign Over[29][18] = 9'b100100100;
assign Over[29][19] = 9'b101101101;
assign Over[29][20] = 9'b110010001;
assign Over[29][21] = 9'b110010001;
assign Over[29][22] = 9'b110010001;
assign Over[29][23] = 9'b110010001;
assign Over[29][24] = 9'b101101001;
assign Over[29][25] = 9'b110001101;
assign Over[29][26] = 9'b110010010;
assign Over[29][27] = 9'b110110010;
assign Over[29][28] = 9'b110010001;
assign Over[29][29] = 9'b101001001;
assign Over[29][30] = 9'b110010001;
assign Over[29][31] = 9'b110010001;
assign Over[29][32] = 9'b101101101;
assign Over[29][35] = 9'b110001101;
assign Over[29][36] = 9'b101101101;
assign Over[29][37] = 9'b100000000;
assign Over[29][38] = 9'b100000000;
assign Over[29][39] = 9'b100000000;
assign Over[29][40] = 9'b100000000;
assign Over[29][41] = 9'b100000000;
assign Over[29][42] = 9'b100100100;
assign Over[29][43] = 9'b110001101;
assign Over[29][44] = 9'b110010001;
assign Over[29][45] = 9'b101101101;
assign Over[29][46] = 9'b110001101;
assign Over[29][47] = 9'b101101101;
assign Over[29][48] = 9'b110010001;
assign Over[29][49] = 9'b110010001;
assign Over[29][50] = 9'b101101101;
assign Over[29][51] = 9'b110010001;
assign Over[29][52] = 9'b101001000;
assign Over[29][53] = 9'b100100100;
assign Over[29][54] = 9'b101101101;
assign Over[29][55] = 9'b101101101;
assign Over[30][15] = 9'b101001001;
assign Over[30][16] = 9'b101101101;
assign Over[30][17] = 9'b100100100;
assign Over[30][18] = 9'b100100100;
assign Over[30][19] = 9'b101101101;
assign Over[30][20] = 9'b110001101;
assign Over[30][21] = 9'b110010001;
assign Over[30][22] = 9'b101101001;
assign Over[30][23] = 9'b110010001;
assign Over[30][24] = 9'b101101101;
assign Over[30][25] = 9'b110010001;
assign Over[30][26] = 9'b101101101;
assign Over[30][27] = 9'b101101101;
assign Over[30][28] = 9'b110010001;
assign Over[30][29] = 9'b101101001;
assign Over[30][30] = 9'b110010001;
assign Over[30][31] = 9'b101101101;
assign Over[30][35] = 9'b110010001;
assign Over[30][36] = 9'b101101101;
assign Over[30][37] = 9'b100000000;
assign Over[30][38] = 9'b100000000;
assign Over[30][39] = 9'b100000000;
assign Over[30][40] = 9'b100000000;
assign Over[30][41] = 9'b100000000;
assign Over[30][42] = 9'b100100100;
assign Over[30][43] = 9'b101101101;
assign Over[30][44] = 9'b110010001;
assign Over[30][45] = 9'b110010001;
assign Over[30][46] = 9'b110010001;
assign Over[30][47] = 9'b101101001;
assign Over[30][48] = 9'b110001101;
assign Over[30][49] = 9'b101101101;
assign Over[30][50] = 9'b101001000;
assign Over[30][51] = 9'b110010001;
assign Over[30][52] = 9'b101001000;
assign Over[30][53] = 9'b100100100;
assign Over[30][54] = 9'b101101101;
assign Over[30][55] = 9'b101101101;
assign Over[31][15] = 9'b101001001;
assign Over[31][16] = 9'b101101101;
assign Over[31][17] = 9'b100100100;
assign Over[31][18] = 9'b100100100;
assign Over[31][19] = 9'b101101101;
assign Over[31][20] = 9'b110001101;
assign Over[31][21] = 9'b110010001;
assign Over[31][22] = 9'b101001001;
assign Over[31][23] = 9'b110010001;
assign Over[31][24] = 9'b101101101;
assign Over[31][25] = 9'b110010001;
assign Over[31][26] = 9'b101001001;
assign Over[31][28] = 9'b110010001;
assign Over[31][29] = 9'b101101101;
assign Over[31][30] = 9'b110010001;
assign Over[31][31] = 9'b101101101;
assign Over[31][35] = 9'b110110010;
assign Over[31][36] = 9'b101101101;
assign Over[31][37] = 9'b100000000;
assign Over[31][38] = 9'b100000000;
assign Over[31][39] = 9'b100000000;
assign Over[31][40] = 9'b100000000;
assign Over[31][41] = 9'b100000000;
assign Over[31][42] = 9'b100100100;
assign Over[31][43] = 9'b101101101;
assign Over[31][44] = 9'b110010001;
assign Over[31][45] = 9'b110010001;
assign Over[31][46] = 9'b110010001;
assign Over[31][47] = 9'b101001001;
assign Over[31][48] = 9'b110001101;
assign Over[31][49] = 9'b101101101;
assign Over[31][50] = 9'b101000100;
assign Over[31][51] = 9'b110010001;
assign Over[31][52] = 9'b101001000;
assign Over[31][53] = 9'b100100100;
assign Over[31][54] = 9'b110001101;
assign Over[31][55] = 9'b101101101;
assign Over[32][15] = 9'b101001001;
assign Over[32][16] = 9'b101101101;
assign Over[32][17] = 9'b100100100;
assign Over[32][18] = 9'b100100100;
assign Over[32][19] = 9'b101101101;
assign Over[32][20] = 9'b110001101;
assign Over[32][21] = 9'b110010001;
assign Over[32][22] = 9'b101001001;
assign Over[32][23] = 9'b110010001;
assign Over[32][24] = 9'b101101101;
assign Over[32][25] = 9'b110010001;
assign Over[32][28] = 9'b110110010;
assign Over[32][29] = 9'b110001101;
assign Over[32][30] = 9'b110010001;
assign Over[32][31] = 9'b110001101;
assign Over[32][36] = 9'b101101101;
assign Over[32][37] = 9'b100000000;
assign Over[32][38] = 9'b100000000;
assign Over[32][39] = 9'b100000000;
assign Over[32][40] = 9'b100000000;
assign Over[32][41] = 9'b100000000;
assign Over[32][42] = 9'b100100100;
assign Over[32][43] = 9'b110001101;
assign Over[32][44] = 9'b101101101;
assign Over[32][45] = 9'b110110010;
assign Over[32][46] = 9'b110010001;
assign Over[32][47] = 9'b101001000;
assign Over[32][48] = 9'b110001101;
assign Over[32][49] = 9'b101101101;
assign Over[32][50] = 9'b101000100;
assign Over[32][51] = 9'b110010001;
assign Over[32][52] = 9'b101001001;
assign Over[32][53] = 9'b101001001;
assign Over[32][54] = 9'b110010001;
assign Over[33][16] = 9'b101101101;
assign Over[33][17] = 9'b101001000;
assign Over[33][18] = 9'b100100100;
assign Over[33][19] = 9'b101101101;
assign Over[33][20] = 9'b110001101;
assign Over[33][21] = 9'b110010001;
assign Over[33][22] = 9'b101001000;
assign Over[33][23] = 9'b110010001;
assign Over[33][24] = 9'b110001101;
assign Over[33][25] = 9'b110010001;
assign Over[33][28] = 9'b110110010;
assign Over[33][29] = 9'b110001101;
assign Over[33][30] = 9'b110010001;
assign Over[33][31] = 9'b101101101;
assign Over[33][36] = 9'b110001101;
assign Over[33][37] = 9'b100100100;
assign Over[33][38] = 9'b100000000;
assign Over[33][39] = 9'b100000000;
assign Over[33][40] = 9'b100000000;
assign Over[33][41] = 9'b100000000;
assign Over[33][42] = 9'b101000100;
assign Over[33][43] = 9'b110010001;
assign Over[33][44] = 9'b101001000;
assign Over[33][45] = 9'b110110110;
assign Over[33][46] = 9'b110010001;
assign Over[33][47] = 9'b100100100;
assign Over[33][48] = 9'b110001101;
assign Over[33][49] = 9'b101101001;
assign Over[33][50] = 9'b100100100;
assign Over[33][51] = 9'b110010001;
assign Over[33][52] = 9'b101101101;
assign Over[33][53] = 9'b110010001;
assign Over[33][54] = 9'b101101101;
assign Over[34][16] = 9'b101101101;
assign Over[34][17] = 9'b110010001;
assign Over[34][18] = 9'b100100100;
assign Over[34][19] = 9'b101101101;
assign Over[34][20] = 9'b101101101;
assign Over[34][21] = 9'b110010001;
assign Over[34][22] = 9'b101001000;
assign Over[34][23] = 9'b110010001;
assign Over[34][24] = 9'b110010001;
assign Over[34][25] = 9'b110010001;
assign Over[34][28] = 9'b110001101;
assign Over[34][29] = 9'b110010001;
assign Over[34][30] = 9'b110010001;
assign Over[34][31] = 9'b101101101;
assign Over[34][36] = 9'b110001101;
assign Over[34][37] = 9'b101101101;
assign Over[34][38] = 9'b100000000;
assign Over[34][39] = 9'b100000000;
assign Over[34][40] = 9'b100000000;
assign Over[34][41] = 9'b100000000;
assign Over[34][42] = 9'b101101101;
assign Over[34][43] = 9'b110010001;
assign Over[34][45] = 9'b110110010;
assign Over[34][46] = 9'b110010001;
assign Over[34][47] = 9'b100000000;
assign Over[34][48] = 9'b110001101;
assign Over[34][49] = 9'b101101001;
assign Over[34][50] = 9'b100100100;
assign Over[34][51] = 9'b110010001;
assign Over[34][52] = 9'b111111111;
assign Over[34][53] = 9'b101101101;
assign Over[35][16] = 9'b100100100;
assign Over[35][17] = 9'b110001101;
assign Over[35][18] = 9'b110010001;
assign Over[35][19] = 9'b110010001;
assign Over[35][20] = 9'b101101101;
assign Over[35][21] = 9'b110010001;
assign Over[35][22] = 9'b101001000;
assign Over[35][23] = 9'b110010001;
assign Over[35][24] = 9'b110010001;
assign Over[35][25] = 9'b110010001;
assign Over[35][29] = 9'b110001101;
assign Over[35][30] = 9'b110010001;
assign Over[35][31] = 9'b101101101;
assign Over[35][36] = 9'b101001001;
assign Over[35][37] = 9'b110010001;
assign Over[35][38] = 9'b101001001;
assign Over[35][39] = 9'b100100100;
assign Over[35][40] = 9'b100100100;
assign Over[35][41] = 9'b101101001;
assign Over[35][42] = 9'b110010001;
assign Over[35][45] = 9'b110010001;
assign Over[35][46] = 9'b101101101;
assign Over[35][48] = 9'b110001101;
assign Over[35][49] = 9'b101101101;
assign Over[35][50] = 9'b101001000;
assign Over[35][51] = 9'b110010001;
assign Over[35][52] = 9'b110010001;
assign Over[35][53] = 9'b110010001;
assign Over[36][17] = 9'b100100100;
assign Over[36][18] = 9'b101101101;
assign Over[36][19] = 9'b110010010;
assign Over[36][20] = 9'b101001001;
assign Over[36][21] = 9'b101101101;
assign Over[36][23] = 9'b101101101;
assign Over[36][24] = 9'b110001101;
assign Over[36][25] = 9'b101101101;
assign Over[36][29] = 9'b101101101;
assign Over[36][30] = 9'b101101101;
assign Over[36][31] = 9'b110110110;
assign Over[36][32] = 9'b101101101;
assign Over[36][37] = 9'b101001001;
assign Over[36][38] = 9'b110010001;
assign Over[36][39] = 9'b110010001;
assign Over[36][40] = 9'b110010001;
assign Over[36][41] = 9'b110001101;
assign Over[36][42] = 9'b101001001;
assign Over[36][45] = 9'b101101101;
assign Over[36][48] = 9'b101101101;
assign Over[36][49] = 9'b110110110;
assign Over[36][50] = 9'b101101101;
assign Over[36][51] = 9'b101101101;
assign Over[36][52] = 9'b101001000;
assign Over[36][53] = 9'b110001101;
assign Over[36][54] = 9'b101101101;
assign Over[37][19] = 9'b101001000;
assign Over[37][30] = 9'b100100100;
assign Over[37][31] = 9'b101001000;
assign Over[37][32] = 9'b100100100;
assign Over[37][38] = 9'b100100100;
assign Over[37][39] = 9'b101001001;
assign Over[37][40] = 9'b101101001;
assign Over[37][49] = 9'b101001000;
assign Over[37][50] = 9'b101001000;
//Total de Lineas = 1053

endmodule
