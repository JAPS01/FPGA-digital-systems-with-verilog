`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:53:22 04/30/2021 
// Design Name: 
// Module Name:    User 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module User(
input enable,
input clock,
input [9:0] X, Y,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg imagen);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= X & hcount < X + RESOLUCION_X & vcount >= Y & vcount < Y + RESOLUCION_Y)
		begin
			if (User[vcount - Y][hcount - X][8] == 1'b1)
			begin
				red   <= User[vcount- Y][hcount- X][7:5];
				green <= User[vcount- Y][hcount- X][4:2];
            blue 	<= User[vcount- Y][hcount- X][1:0];
				imagen  <= 1'b1;
			end
			else
				imagen <= 0;
			end
		else
		imagen <= 0;
	end
end

parameter RESOLUCION_X = 72;
parameter RESOLUCION_Y = 25;
wire [8:0] User[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign User[0][0] = 9'b111111111;
assign User[0][1] = 9'b111111111;
assign User[0][2] = 9'b111111111;
assign User[0][3] = 9'b111111111;
assign User[0][4] = 9'b111111111;
assign User[0][5] = 9'b111111111;
assign User[0][6] = 9'b111111111;
assign User[0][7] = 9'b111111111;
assign User[0][8] = 9'b111111111;
assign User[0][9] = 9'b111111111;
assign User[0][10] = 9'b111111111;
assign User[0][11] = 9'b111111111;
assign User[0][12] = 9'b111111111;
assign User[0][13] = 9'b111111111;
assign User[0][14] = 9'b111111111;
assign User[0][15] = 9'b111111111;
assign User[0][16] = 9'b111111111;
assign User[0][17] = 9'b111111111;
assign User[0][18] = 9'b111111111;
assign User[0][19] = 9'b111111111;
assign User[0][20] = 9'b111111111;
assign User[0][21] = 9'b111111111;
assign User[0][22] = 9'b111111111;
assign User[0][23] = 9'b111111111;
assign User[0][24] = 9'b111111111;
assign User[0][25] = 9'b111111111;
assign User[0][26] = 9'b111111111;
assign User[0][27] = 9'b111111111;
assign User[0][28] = 9'b111111111;
assign User[0][29] = 9'b111111111;
assign User[0][30] = 9'b111111111;
assign User[0][31] = 9'b111111111;
assign User[0][32] = 9'b111111111;
assign User[0][33] = 9'b111111111;
assign User[0][34] = 9'b111111111;
assign User[0][35] = 9'b111111111;
assign User[0][36] = 9'b111111111;
assign User[0][37] = 9'b111111111;
assign User[0][38] = 9'b111111111;
assign User[0][39] = 9'b111111111;
assign User[0][40] = 9'b111111111;
assign User[0][41] = 9'b111111111;
assign User[0][42] = 9'b111111111;
assign User[0][43] = 9'b111111111;
assign User[0][44] = 9'b111111111;
assign User[0][45] = 9'b111111111;
assign User[0][46] = 9'b111111111;
assign User[0][47] = 9'b111111111;
assign User[0][48] = 9'b111111111;
assign User[0][49] = 9'b111111111;
assign User[0][50] = 9'b111111111;
assign User[0][51] = 9'b111111111;
assign User[0][52] = 9'b111111111;
assign User[0][53] = 9'b111111111;
assign User[0][54] = 9'b111111111;
assign User[0][55] = 9'b111111111;
assign User[0][56] = 9'b111111111;
assign User[0][57] = 9'b111111111;
assign User[0][58] = 9'b111111111;
assign User[0][59] = 9'b111111111;
assign User[0][60] = 9'b111111111;
assign User[0][61] = 9'b111111111;
assign User[0][62] = 9'b111111111;
assign User[0][63] = 9'b111111111;
assign User[0][64] = 9'b111111111;
assign User[0][65] = 9'b111111111;
assign User[0][66] = 9'b111111111;
assign User[0][67] = 9'b111111111;
assign User[0][68] = 9'b111111111;
assign User[0][69] = 9'b111111111;
assign User[0][70] = 9'b111111111;
assign User[0][71] = 9'b111111111;
assign User[1][0] = 9'b111111111;
assign User[1][1] = 9'b111111111;
assign User[1][2] = 9'b111111111;
assign User[1][3] = 9'b111111111;
assign User[1][4] = 9'b111111111;
assign User[1][5] = 9'b111111111;
assign User[1][6] = 9'b111111111;
assign User[1][7] = 9'b111111111;
assign User[1][8] = 9'b111111111;
assign User[1][9] = 9'b111111111;
assign User[1][10] = 9'b111111111;
assign User[1][11] = 9'b111111111;
assign User[1][12] = 9'b111111111;
assign User[1][13] = 9'b111111111;
assign User[1][14] = 9'b111111111;
assign User[1][15] = 9'b111111111;
assign User[1][16] = 9'b111111111;
assign User[1][17] = 9'b111111111;
assign User[1][18] = 9'b111111111;
assign User[1][19] = 9'b111111111;
assign User[1][20] = 9'b111111111;
assign User[1][21] = 9'b111111111;
assign User[1][22] = 9'b111111111;
assign User[1][23] = 9'b111111111;
assign User[1][24] = 9'b111111111;
assign User[1][25] = 9'b111111111;
assign User[1][26] = 9'b111111111;
assign User[1][27] = 9'b111111111;
assign User[1][28] = 9'b111111111;
assign User[1][29] = 9'b111111111;
assign User[1][30] = 9'b111111111;
assign User[1][31] = 9'b111111111;
assign User[1][32] = 9'b111111111;
assign User[1][33] = 9'b111111111;
assign User[1][34] = 9'b111111111;
assign User[1][35] = 9'b111111111;
assign User[1][36] = 9'b111111111;
assign User[1][37] = 9'b111111111;
assign User[1][38] = 9'b111111111;
assign User[1][39] = 9'b111111111;
assign User[1][40] = 9'b111111111;
assign User[1][41] = 9'b111111111;
assign User[1][42] = 9'b111111111;
assign User[1][43] = 9'b111111111;
assign User[1][44] = 9'b111111111;
assign User[1][45] = 9'b111111111;
assign User[1][46] = 9'b111111111;
assign User[1][47] = 9'b111111111;
assign User[1][48] = 9'b111111111;
assign User[1][49] = 9'b111111111;
assign User[1][50] = 9'b111111111;
assign User[1][51] = 9'b111111111;
assign User[1][52] = 9'b111111111;
assign User[1][53] = 9'b111111111;
assign User[1][54] = 9'b111111111;
assign User[1][55] = 9'b111111111;
assign User[1][56] = 9'b111111111;
assign User[1][57] = 9'b111111111;
assign User[1][58] = 9'b111111111;
assign User[1][59] = 9'b111111111;
assign User[1][60] = 9'b111111111;
assign User[1][61] = 9'b111111111;
assign User[1][62] = 9'b111111111;
assign User[1][63] = 9'b111111111;
assign User[1][64] = 9'b111111111;
assign User[1][65] = 9'b111111111;
assign User[1][66] = 9'b111111111;
assign User[1][67] = 9'b111111111;
assign User[1][68] = 9'b111111111;
assign User[1][69] = 9'b111111111;
assign User[1][70] = 9'b111111111;
assign User[1][71] = 9'b111111111;
assign User[2][0] = 9'b111111111;
assign User[2][1] = 9'b111111111;
assign User[2][2] = 9'b111111111;
assign User[2][3] = 9'b111111111;
assign User[2][4] = 9'b111111111;
assign User[2][5] = 9'b111111111;
assign User[2][6] = 9'b111111111;
assign User[2][7] = 9'b111111111;
assign User[2][8] = 9'b111111111;
assign User[2][9] = 9'b111111111;
assign User[2][10] = 9'b111111111;
assign User[2][11] = 9'b111111111;
assign User[2][12] = 9'b111111111;
assign User[2][13] = 9'b111111111;
assign User[2][14] = 9'b111111111;
assign User[2][15] = 9'b111111111;
assign User[2][16] = 9'b111111111;
assign User[2][17] = 9'b111111111;
assign User[2][18] = 9'b111111111;
assign User[2][19] = 9'b111111111;
assign User[2][20] = 9'b111111111;
assign User[2][21] = 9'b111111111;
assign User[2][22] = 9'b111111111;
assign User[2][23] = 9'b111111111;
assign User[2][24] = 9'b111111111;
assign User[2][25] = 9'b111111111;
assign User[2][26] = 9'b111111111;
assign User[2][27] = 9'b111111111;
assign User[2][28] = 9'b111111111;
assign User[2][29] = 9'b111111111;
assign User[2][30] = 9'b111111111;
assign User[2][31] = 9'b111111111;
assign User[2][32] = 9'b111111111;
assign User[2][33] = 9'b111111111;
assign User[2][34] = 9'b111111111;
assign User[2][35] = 9'b111111111;
assign User[2][36] = 9'b111111111;
assign User[2][37] = 9'b111111111;
assign User[2][38] = 9'b111111111;
assign User[2][39] = 9'b111111111;
assign User[2][40] = 9'b111111111;
assign User[2][41] = 9'b111111111;
assign User[2][42] = 9'b111111111;
assign User[2][43] = 9'b111111111;
assign User[2][44] = 9'b111111111;
assign User[2][45] = 9'b111111111;
assign User[2][46] = 9'b111111111;
assign User[2][47] = 9'b111111111;
assign User[2][48] = 9'b111111111;
assign User[2][49] = 9'b111111111;
assign User[2][50] = 9'b111111111;
assign User[2][51] = 9'b111111111;
assign User[2][52] = 9'b111111111;
assign User[2][53] = 9'b111111111;
assign User[2][54] = 9'b111111111;
assign User[2][55] = 9'b111111111;
assign User[2][56] = 9'b111111111;
assign User[2][57] = 9'b111111111;
assign User[2][58] = 9'b111111111;
assign User[2][59] = 9'b111111111;
assign User[2][60] = 9'b111111111;
assign User[2][61] = 9'b111111111;
assign User[2][62] = 9'b111111111;
assign User[2][63] = 9'b111111111;
assign User[2][64] = 9'b111111111;
assign User[2][65] = 9'b111111111;
assign User[2][66] = 9'b111111111;
assign User[2][67] = 9'b111111111;
assign User[2][68] = 9'b111111111;
assign User[2][69] = 9'b111111111;
assign User[2][70] = 9'b111111111;
assign User[2][71] = 9'b111111111;
assign User[3][0] = 9'b111111111;
assign User[3][1] = 9'b111111111;
assign User[3][2] = 9'b111111111;
assign User[3][3] = 9'b111111111;
assign User[3][4] = 9'b111111111;
assign User[3][5] = 9'b111111111;
assign User[3][6] = 9'b111111111;
assign User[3][7] = 9'b111111111;
assign User[3][8] = 9'b111111111;
assign User[3][9] = 9'b111111111;
assign User[3][10] = 9'b111111111;
assign User[3][11] = 9'b111111111;
assign User[3][12] = 9'b111111111;
assign User[3][13] = 9'b111111111;
assign User[3][14] = 9'b111111111;
assign User[3][15] = 9'b111111111;
assign User[3][16] = 9'b111111111;
assign User[3][17] = 9'b111111111;
assign User[3][18] = 9'b111111111;
assign User[3][19] = 9'b101101101;
assign User[3][20] = 9'b101001001;
assign User[3][21] = 9'b111111111;
assign User[3][22] = 9'b111111111;
assign User[3][23] = 9'b111111111;
assign User[3][24] = 9'b111111111;
assign User[3][25] = 9'b111111111;
assign User[3][26] = 9'b111111111;
assign User[3][27] = 9'b111111111;
assign User[3][28] = 9'b111111111;
assign User[3][29] = 9'b111111111;
assign User[3][30] = 9'b111111111;
assign User[3][31] = 9'b111111111;
assign User[3][32] = 9'b111111111;
assign User[3][33] = 9'b111111111;
assign User[3][34] = 9'b111111111;
assign User[3][35] = 9'b111111111;
assign User[3][36] = 9'b111111111;
assign User[3][37] = 9'b111111111;
assign User[3][38] = 9'b111111111;
assign User[3][39] = 9'b111111111;
assign User[3][40] = 9'b111111111;
assign User[3][41] = 9'b111111111;
assign User[3][42] = 9'b111111111;
assign User[3][43] = 9'b111111111;
assign User[3][44] = 9'b111111111;
assign User[3][45] = 9'b111111111;
assign User[3][46] = 9'b111111111;
assign User[3][47] = 9'b111111111;
assign User[3][48] = 9'b111111111;
assign User[3][49] = 9'b111111111;
assign User[3][50] = 9'b111111111;
assign User[3][51] = 9'b111111111;
assign User[3][52] = 9'b111111111;
assign User[3][53] = 9'b111111111;
assign User[3][54] = 9'b111111111;
assign User[3][55] = 9'b111111111;
assign User[3][56] = 9'b111111111;
assign User[3][57] = 9'b111111111;
assign User[3][58] = 9'b111111111;
assign User[3][59] = 9'b111111111;
assign User[3][60] = 9'b111111111;
assign User[3][61] = 9'b111111111;
assign User[3][62] = 9'b111111111;
assign User[3][63] = 9'b111111111;
assign User[3][64] = 9'b111111111;
assign User[3][65] = 9'b111111111;
assign User[3][66] = 9'b111111111;
assign User[3][67] = 9'b111111111;
assign User[3][68] = 9'b111111111;
assign User[3][69] = 9'b111111111;
assign User[3][70] = 9'b111111111;
assign User[3][71] = 9'b111111111;
assign User[4][0] = 9'b111111111;
assign User[4][1] = 9'b111111111;
assign User[4][2] = 9'b111111111;
assign User[4][3] = 9'b111111111;
assign User[4][4] = 9'b111111111;
assign User[4][5] = 9'b101101101;
assign User[4][6] = 9'b100100100;
assign User[4][7] = 9'b111111111;
assign User[4][8] = 9'b101001001;
assign User[4][9] = 9'b101101101;
assign User[4][10] = 9'b111111111;
assign User[4][11] = 9'b101001000;
assign User[4][12] = 9'b100100100;
assign User[4][13] = 9'b100100100;
assign User[4][14] = 9'b101001001;
assign User[4][15] = 9'b110010001;
assign User[4][16] = 9'b100100100;
assign User[4][17] = 9'b110110110;
assign User[4][18] = 9'b111111111;
assign User[4][19] = 9'b101101101;
assign User[4][20] = 9'b110010001;
assign User[4][21] = 9'b100100100;
assign User[4][22] = 9'b101101101;
assign User[4][23] = 9'b101101101;
assign User[4][24] = 9'b100000000;
assign User[4][25] = 9'b110010001;
assign User[4][26] = 9'b101101101;
assign User[4][27] = 9'b101101101;
assign User[4][28] = 9'b111111111;
assign User[4][29] = 9'b111111111;
assign User[4][30] = 9'b111111111;
assign User[4][31] = 9'b110010010;
assign User[4][32] = 9'b100100100;
assign User[4][33] = 9'b110010010;
assign User[4][34] = 9'b111111111;
assign User[4][35] = 9'b111111111;
assign User[4][36] = 9'b111111111;
assign User[4][37] = 9'b111111111;
assign User[4][38] = 9'b111111111;
assign User[4][39] = 9'b111111111;
assign User[4][40] = 9'b110010001;
assign User[4][41] = 9'b101001001;
assign User[4][42] = 9'b101101101;
assign User[4][43] = 9'b101001001;
assign User[4][44] = 9'b101101101;
assign User[4][45] = 9'b100100100;
assign User[4][46] = 9'b100100100;
assign User[4][47] = 9'b100100100;
assign User[4][48] = 9'b110010010;
assign User[4][49] = 9'b101101101;
assign User[4][50] = 9'b100100100;
assign User[4][51] = 9'b111111111;
assign User[4][52] = 9'b111111111;
assign User[4][53] = 9'b110010010;
assign User[4][54] = 9'b100000000;
assign User[4][55] = 9'b110110110;
assign User[4][56] = 9'b111111111;
assign User[4][57] = 9'b110010010;
assign User[4][58] = 9'b100100100;
assign User[4][59] = 9'b110010010;
assign User[4][60] = 9'b111111111;
assign User[4][61] = 9'b111111111;
assign User[4][62] = 9'b110010001;
assign User[4][63] = 9'b101001001;
assign User[4][64] = 9'b101101101;
assign User[4][65] = 9'b101001000;
assign User[4][66] = 9'b111111111;
assign User[4][67] = 9'b111111111;
assign User[4][68] = 9'b111111111;
assign User[4][69] = 9'b111111111;
assign User[4][70] = 9'b111111111;
assign User[4][71] = 9'b111111111;
assign User[5][0] = 9'b111111111;
assign User[5][1] = 9'b111111111;
assign User[5][2] = 9'b111111111;
assign User[5][3] = 9'b111111111;
assign User[5][4] = 9'b111111111;
assign User[5][5] = 9'b110010010;
assign User[5][6] = 9'b101001001;
assign User[5][7] = 9'b111111111;
assign User[5][8] = 9'b110010001;
assign User[5][9] = 9'b111111111;
assign User[5][10] = 9'b111111111;
assign User[5][11] = 9'b101001001;
assign User[5][12] = 9'b101101101;
assign User[5][13] = 9'b110110110;
assign User[5][14] = 9'b110110110;
assign User[5][15] = 9'b111111111;
assign User[5][16] = 9'b101001001;
assign User[5][17] = 9'b110110110;
assign User[5][18] = 9'b111111111;
assign User[5][19] = 9'b110010001;
assign User[5][20] = 9'b111111111;
assign User[5][21] = 9'b100100100;
assign User[5][22] = 9'b110010010;
assign User[5][23] = 9'b110110110;
assign User[5][24] = 9'b100100100;
assign User[5][25] = 9'b101101101;
assign User[5][26] = 9'b110110110;
assign User[5][27] = 9'b110110110;
assign User[5][28] = 9'b111111111;
assign User[5][29] = 9'b111111111;
assign User[5][30] = 9'b111111111;
assign User[5][31] = 9'b110010010;
assign User[5][32] = 9'b100100100;
assign User[5][33] = 9'b110010001;
assign User[5][34] = 9'b111111111;
assign User[5][35] = 9'b111111111;
assign User[5][36] = 9'b111111111;
assign User[5][37] = 9'b111111111;
assign User[5][38] = 9'b111111111;
assign User[5][39] = 9'b111111111;
assign User[5][40] = 9'b101001001;
assign User[5][41] = 9'b110010001;
assign User[5][42] = 9'b111111111;
assign User[5][43] = 9'b110110110;
assign User[5][44] = 9'b111111111;
assign User[5][45] = 9'b101001000;
assign User[5][46] = 9'b111111111;
assign User[5][47] = 9'b110010010;
assign User[5][48] = 9'b111111111;
assign User[5][49] = 9'b110010010;
assign User[5][50] = 9'b100100100;
assign User[5][51] = 9'b111111111;
assign User[5][52] = 9'b111111111;
assign User[5][53] = 9'b111111111;
assign User[5][54] = 9'b100000000;
assign User[5][55] = 9'b111111111;
assign User[5][56] = 9'b111111111;
assign User[5][57] = 9'b110010010;
assign User[5][58] = 9'b100100100;
assign User[5][59] = 9'b110010001;
assign User[5][60] = 9'b111111111;
assign User[5][61] = 9'b111111111;
assign User[5][62] = 9'b101001001;
assign User[5][63] = 9'b110010001;
assign User[5][64] = 9'b111111111;
assign User[5][65] = 9'b110110110;
assign User[5][66] = 9'b111111111;
assign User[5][67] = 9'b111111111;
assign User[5][68] = 9'b111111111;
assign User[5][69] = 9'b111111111;
assign User[5][70] = 9'b111111111;
assign User[5][71] = 9'b111111111;
assign User[6][0] = 9'b111111111;
assign User[6][1] = 9'b111111111;
assign User[6][2] = 9'b111111111;
assign User[6][3] = 9'b111111111;
assign User[6][4] = 9'b111111111;
assign User[6][5] = 9'b110010010;
assign User[6][6] = 9'b101001000;
assign User[6][7] = 9'b100100100;
assign User[6][8] = 9'b101101101;
assign User[6][9] = 9'b111111111;
assign User[6][10] = 9'b111111111;
assign User[6][11] = 9'b100100100;
assign User[6][12] = 9'b101001000;
assign User[6][13] = 9'b101001000;
assign User[6][14] = 9'b111111111;
assign User[6][15] = 9'b111111111;
assign User[6][16] = 9'b110010001;
assign User[6][17] = 9'b101101101;
assign User[6][18] = 9'b110110110;
assign User[6][19] = 9'b110110110;
assign User[6][20] = 9'b111111111;
assign User[6][21] = 9'b100100100;
assign User[6][22] = 9'b110010010;
assign User[6][23] = 9'b110110110;
assign User[6][24] = 9'b110010001;
assign User[6][25] = 9'b100100100;
assign User[6][26] = 9'b101101101;
assign User[6][27] = 9'b111111111;
assign User[6][28] = 9'b111111111;
assign User[6][29] = 9'b111111111;
assign User[6][30] = 9'b110110110;
assign User[6][31] = 9'b101001000;
assign User[6][32] = 9'b101101101;
assign User[6][33] = 9'b100100100;
assign User[6][34] = 9'b110010001;
assign User[6][35] = 9'b111111111;
assign User[6][36] = 9'b111111111;
assign User[6][37] = 9'b111111111;
assign User[6][38] = 9'b111111111;
assign User[6][39] = 9'b111111111;
assign User[6][40] = 9'b110010010;
assign User[6][41] = 9'b100100100;
assign User[6][42] = 9'b101101101;
assign User[6][43] = 9'b110110110;
assign User[6][44] = 9'b101101101;
assign User[6][45] = 9'b100100100;
assign User[6][46] = 9'b101001000;
assign User[6][47] = 9'b110010001;
assign User[6][48] = 9'b111111111;
assign User[6][49] = 9'b110010001;
assign User[6][50] = 9'b100100100;
assign User[6][51] = 9'b111111111;
assign User[6][52] = 9'b111111111;
assign User[6][53] = 9'b111111111;
assign User[6][54] = 9'b100000000;
assign User[6][55] = 9'b111111111;
assign User[6][56] = 9'b110110110;
assign User[6][57] = 9'b101001000;
assign User[6][58] = 9'b101101101;
assign User[6][59] = 9'b100100100;
assign User[6][60] = 9'b110010001;
assign User[6][61] = 9'b111111111;
assign User[6][62] = 9'b110010010;
assign User[6][63] = 9'b100100100;
assign User[6][64] = 9'b101101101;
assign User[6][65] = 9'b110110110;
assign User[6][66] = 9'b111111111;
assign User[6][67] = 9'b111111111;
assign User[6][68] = 9'b111111111;
assign User[6][69] = 9'b111111111;
assign User[6][70] = 9'b111111111;
assign User[6][71] = 9'b111111111;
assign User[7][0] = 9'b111111111;
assign User[7][1] = 9'b111111111;
assign User[7][2] = 9'b111111111;
assign User[7][3] = 9'b111111111;
assign User[7][4] = 9'b111111111;
assign User[7][5] = 9'b110010010;
assign User[7][6] = 9'b101001000;
assign User[7][7] = 9'b110010001;
assign User[7][8] = 9'b100100100;
assign User[7][9] = 9'b111111111;
assign User[7][10] = 9'b111111111;
assign User[7][11] = 9'b100100100;
assign User[7][12] = 9'b101001001;
assign User[7][13] = 9'b110010001;
assign User[7][14] = 9'b111111111;
assign User[7][15] = 9'b111111111;
assign User[7][16] = 9'b111111111;
assign User[7][17] = 9'b101001000;
assign User[7][18] = 9'b101101101;
assign User[7][19] = 9'b111111111;
assign User[7][20] = 9'b111111111;
assign User[7][21] = 9'b101001000;
assign User[7][22] = 9'b110010010;
assign User[7][23] = 9'b110110110;
assign User[7][24] = 9'b111111111;
assign User[7][25] = 9'b101101101;
assign User[7][26] = 9'b100100100;
assign User[7][27] = 9'b111111111;
assign User[7][28] = 9'b111111111;
assign User[7][29] = 9'b111111111;
assign User[7][30] = 9'b111111111;
assign User[7][31] = 9'b101101101;
assign User[7][32] = 9'b101001000;
assign User[7][33] = 9'b100100100;
assign User[7][34] = 9'b110010001;
assign User[7][35] = 9'b111111111;
assign User[7][36] = 9'b111111111;
assign User[7][37] = 9'b111111111;
assign User[7][38] = 9'b111111111;
assign User[7][39] = 9'b111111111;
assign User[7][40] = 9'b111111111;
assign User[7][41] = 9'b110110110;
assign User[7][42] = 9'b101101101;
assign User[7][43] = 9'b100100100;
assign User[7][44] = 9'b100100100;
assign User[7][45] = 9'b100100100;
assign User[7][46] = 9'b101101101;
assign User[7][47] = 9'b111111111;
assign User[7][48] = 9'b111111111;
assign User[7][49] = 9'b110010010;
assign User[7][50] = 9'b101001000;
assign User[7][51] = 9'b110110110;
assign User[7][52] = 9'b101101101;
assign User[7][53] = 9'b111111111;
assign User[7][54] = 9'b100100100;
assign User[7][55] = 9'b111111111;
assign User[7][56] = 9'b111111111;
assign User[7][57] = 9'b101101101;
assign User[7][58] = 9'b101001000;
assign User[7][59] = 9'b100100100;
assign User[7][60] = 9'b110010001;
assign User[7][61] = 9'b111111111;
assign User[7][62] = 9'b111111111;
assign User[7][63] = 9'b110110110;
assign User[7][64] = 9'b101101101;
assign User[7][65] = 9'b100100100;
assign User[7][66] = 9'b110110110;
assign User[7][67] = 9'b111111111;
assign User[7][68] = 9'b111111111;
assign User[7][69] = 9'b111111111;
assign User[7][70] = 9'b111111111;
assign User[7][71] = 9'b111111111;
assign User[8][0] = 9'b111111111;
assign User[8][1] = 9'b111111111;
assign User[8][2] = 9'b111111111;
assign User[8][3] = 9'b111111111;
assign User[8][4] = 9'b111111111;
assign User[8][5] = 9'b101101101;
assign User[8][6] = 9'b100100100;
assign User[8][7] = 9'b111111111;
assign User[8][8] = 9'b100100100;
assign User[8][9] = 9'b101001000;
assign User[8][10] = 9'b111111111;
assign User[8][11] = 9'b100100100;
assign User[8][12] = 9'b100100100;
assign User[8][13] = 9'b101101101;
assign User[8][14] = 9'b100100100;
assign User[8][15] = 9'b110110110;
assign User[8][16] = 9'b111111111;
assign User[8][17] = 9'b100100100;
assign User[8][18] = 9'b101001001;
assign User[8][19] = 9'b111111111;
assign User[8][20] = 9'b111111111;
assign User[8][21] = 9'b100000000;
assign User[8][22] = 9'b101101101;
assign User[8][23] = 9'b101101101;
assign User[8][24] = 9'b101101101;
assign User[8][25] = 9'b111111111;
assign User[8][26] = 9'b100100100;
assign User[8][27] = 9'b110110110;
assign User[8][28] = 9'b111111111;
assign User[8][29] = 9'b111111111;
assign User[8][30] = 9'b100100100;
assign User[8][31] = 9'b110010001;
assign User[8][32] = 9'b111111111;
assign User[8][33] = 9'b101001000;
assign User[8][34] = 9'b100100100;
assign User[8][35] = 9'b110110110;
assign User[8][36] = 9'b100100100;
assign User[8][37] = 9'b111111111;
assign User[8][38] = 9'b111111111;
assign User[8][39] = 9'b111111111;
assign User[8][40] = 9'b101001000;
assign User[8][41] = 9'b101101101;
assign User[8][42] = 9'b111111111;
assign User[8][43] = 9'b101001000;
assign User[8][44] = 9'b101001001;
assign User[8][45] = 9'b100000000;
assign User[8][46] = 9'b101101101;
assign User[8][47] = 9'b101001001;
assign User[8][48] = 9'b101001001;
assign User[8][49] = 9'b101101101;
assign User[8][50] = 9'b100100100;
assign User[8][51] = 9'b101101101;
assign User[8][52] = 9'b100100100;
assign User[8][53] = 9'b110010001;
assign User[8][54] = 9'b100100100;
assign User[8][55] = 9'b110110110;
assign User[8][56] = 9'b100100100;
assign User[8][57] = 9'b110010001;
assign User[8][58] = 9'b111111111;
assign User[8][59] = 9'b101001000;
assign User[8][60] = 9'b100100100;
assign User[8][61] = 9'b111111111;
assign User[8][62] = 9'b101001001;
assign User[8][63] = 9'b101101101;
assign User[8][64] = 9'b111111111;
assign User[8][65] = 9'b100100100;
assign User[8][66] = 9'b110110110;
assign User[8][67] = 9'b111111111;
assign User[8][68] = 9'b111111111;
assign User[8][69] = 9'b111111111;
assign User[8][70] = 9'b111111111;
assign User[8][71] = 9'b111111111;
assign User[9][0] = 9'b111111111;
assign User[9][1] = 9'b111111111;
assign User[9][2] = 9'b111111111;
assign User[9][3] = 9'b111111111;
assign User[9][4] = 9'b111111111;
assign User[9][5] = 9'b110010001;
assign User[9][6] = 9'b101101101;
assign User[9][7] = 9'b110110110;
assign User[9][8] = 9'b110010001;
assign User[9][9] = 9'b101101101;
assign User[9][10] = 9'b110010001;
assign User[9][11] = 9'b101101101;
assign User[9][12] = 9'b101101101;
assign User[9][13] = 9'b101101101;
assign User[9][14] = 9'b101101101;
assign User[9][15] = 9'b110110110;
assign User[9][16] = 9'b111111111;
assign User[9][17] = 9'b101101101;
assign User[9][18] = 9'b110010001;
assign User[9][19] = 9'b111111111;
assign User[9][20] = 9'b111111111;
assign User[9][21] = 9'b101101101;
assign User[9][22] = 9'b101101101;
assign User[9][23] = 9'b101101101;
assign User[9][24] = 9'b101101101;
assign User[9][25] = 9'b111111111;
assign User[9][26] = 9'b110010001;
assign User[9][27] = 9'b111111111;
assign User[9][28] = 9'b111111111;
assign User[9][29] = 9'b110110110;
assign User[9][30] = 9'b101101101;
assign User[9][31] = 9'b110010001;
assign User[9][32] = 9'b111111111;
assign User[9][33] = 9'b101101101;
assign User[9][34] = 9'b101101101;
assign User[9][35] = 9'b110010010;
assign User[9][36] = 9'b110010001;
assign User[9][37] = 9'b111111111;
assign User[9][38] = 9'b111111111;
assign User[9][39] = 9'b111111111;
assign User[9][40] = 9'b101101101;
assign User[9][41] = 9'b101101101;
assign User[9][42] = 9'b110010001;
assign User[9][43] = 9'b110110110;
assign User[9][44] = 9'b110010010;
assign User[9][45] = 9'b101101101;
assign User[9][46] = 9'b101101101;
assign User[9][47] = 9'b101101101;
assign User[9][48] = 9'b101101101;
assign User[9][49] = 9'b110010001;
assign User[9][50] = 9'b101101101;
assign User[9][51] = 9'b111111111;
assign User[9][52] = 9'b110010001;
assign User[9][53] = 9'b101101101;
assign User[9][54] = 9'b110110110;
assign User[9][55] = 9'b111111111;
assign User[9][56] = 9'b101101101;
assign User[9][57] = 9'b110010001;
assign User[9][58] = 9'b111111111;
assign User[9][59] = 9'b101101101;
assign User[9][60] = 9'b101101101;
assign User[9][61] = 9'b110010010;
assign User[9][62] = 9'b101101101;
assign User[9][63] = 9'b101101101;
assign User[9][64] = 9'b110010001;
assign User[9][65] = 9'b110110110;
assign User[9][66] = 9'b111111111;
assign User[9][67] = 9'b111111111;
assign User[9][68] = 9'b111111111;
assign User[9][69] = 9'b111111111;
assign User[9][70] = 9'b111111111;
assign User[9][71] = 9'b111111111;
assign User[10][0] = 9'b111111111;
assign User[10][1] = 9'b111111111;
assign User[10][2] = 9'b111111111;
assign User[10][3] = 9'b111111111;
assign User[10][4] = 9'b111111111;
assign User[10][5] = 9'b111111111;
assign User[10][6] = 9'b111111111;
assign User[10][7] = 9'b111111111;
assign User[10][8] = 9'b111111111;
assign User[10][9] = 9'b111111111;
assign User[10][10] = 9'b111111111;
assign User[10][11] = 9'b111111111;
assign User[10][12] = 9'b111111111;
assign User[10][13] = 9'b111111111;
assign User[10][14] = 9'b111111111;
assign User[10][15] = 9'b111111111;
assign User[10][16] = 9'b111111111;
assign User[10][17] = 9'b111111111;
assign User[10][18] = 9'b111111111;
assign User[10][19] = 9'b111111111;
assign User[10][20] = 9'b111111111;
assign User[10][21] = 9'b111111111;
assign User[10][22] = 9'b111111111;
assign User[10][23] = 9'b111111111;
assign User[10][24] = 9'b111111111;
assign User[10][25] = 9'b111111111;
assign User[10][26] = 9'b111111111;
assign User[10][27] = 9'b111111111;
assign User[10][28] = 9'b111111111;
assign User[10][29] = 9'b111111111;
assign User[10][30] = 9'b111111111;
assign User[10][31] = 9'b111111111;
assign User[10][32] = 9'b111111111;
assign User[10][33] = 9'b111111111;
assign User[10][34] = 9'b111111111;
assign User[10][35] = 9'b111111111;
assign User[10][36] = 9'b111111111;
assign User[10][37] = 9'b111111111;
assign User[10][38] = 9'b111111111;
assign User[10][39] = 9'b111111111;
assign User[10][40] = 9'b111111111;
assign User[10][41] = 9'b111111111;
assign User[10][42] = 9'b111111111;
assign User[10][43] = 9'b111111111;
assign User[10][44] = 9'b111111111;
assign User[10][45] = 9'b111111111;
assign User[10][46] = 9'b111111111;
assign User[10][47] = 9'b111111111;
assign User[10][48] = 9'b111111111;
assign User[10][49] = 9'b111111111;
assign User[10][50] = 9'b111111111;
assign User[10][51] = 9'b111111111;
assign User[10][52] = 9'b111111111;
assign User[10][53] = 9'b111111111;
assign User[10][54] = 9'b111111111;
assign User[10][55] = 9'b111111111;
assign User[10][56] = 9'b111111111;
assign User[10][57] = 9'b111111111;
assign User[10][58] = 9'b111111111;
assign User[10][59] = 9'b111111111;
assign User[10][60] = 9'b111111111;
assign User[10][61] = 9'b111111111;
assign User[10][62] = 9'b111111111;
assign User[10][63] = 9'b111111111;
assign User[10][64] = 9'b111111111;
assign User[10][65] = 9'b111111111;
assign User[10][66] = 9'b111111111;
assign User[10][67] = 9'b111111111;
assign User[10][68] = 9'b111111111;
assign User[10][69] = 9'b111111111;
assign User[10][70] = 9'b111111111;
assign User[10][71] = 9'b111111111;
assign User[11][0] = 9'b111111111;
assign User[11][1] = 9'b111111111;
assign User[11][2] = 9'b111111111;
assign User[11][3] = 9'b111111111;
assign User[11][4] = 9'b111111111;
assign User[11][5] = 9'b111111111;
assign User[11][6] = 9'b111111111;
assign User[11][7] = 9'b111111111;
assign User[11][8] = 9'b111111111;
assign User[11][9] = 9'b111111111;
assign User[11][10] = 9'b111111111;
assign User[11][11] = 9'b111111111;
assign User[11][12] = 9'b111111111;
assign User[11][13] = 9'b111111111;
assign User[11][14] = 9'b111111111;
assign User[11][15] = 9'b111111111;
assign User[11][16] = 9'b111111111;
assign User[11][17] = 9'b111111111;
assign User[11][18] = 9'b111111111;
assign User[11][19] = 9'b111111111;
assign User[11][20] = 9'b111111111;
assign User[11][21] = 9'b111111111;
assign User[11][22] = 9'b111111111;
assign User[11][23] = 9'b111111111;
assign User[11][24] = 9'b111111111;
assign User[11][25] = 9'b111111111;
assign User[11][26] = 9'b111111111;
assign User[11][27] = 9'b111111111;
assign User[11][28] = 9'b111111111;
assign User[11][29] = 9'b111111111;
assign User[11][30] = 9'b111111111;
assign User[11][31] = 9'b111111111;
assign User[11][32] = 9'b111111111;
assign User[11][33] = 9'b111111111;
assign User[11][34] = 9'b111111111;
assign User[11][35] = 9'b111111111;
assign User[11][36] = 9'b111111111;
assign User[11][37] = 9'b111111111;
assign User[11][38] = 9'b111111111;
assign User[11][39] = 9'b111111111;
assign User[11][40] = 9'b111111111;
assign User[11][41] = 9'b111111111;
assign User[11][42] = 9'b111111111;
assign User[11][43] = 9'b111111111;
assign User[11][44] = 9'b111111111;
assign User[11][45] = 9'b111111111;
assign User[11][46] = 9'b111111111;
assign User[11][47] = 9'b111111111;
assign User[11][48] = 9'b111111111;
assign User[11][49] = 9'b111111111;
assign User[11][50] = 9'b111111111;
assign User[11][51] = 9'b111111111;
assign User[11][52] = 9'b111111111;
assign User[11][53] = 9'b111111111;
assign User[11][54] = 9'b111111111;
assign User[11][55] = 9'b111111111;
assign User[11][56] = 9'b111111111;
assign User[11][57] = 9'b111111111;
assign User[11][58] = 9'b111111111;
assign User[11][59] = 9'b111111111;
assign User[11][60] = 9'b111111111;
assign User[11][61] = 9'b111111111;
assign User[11][62] = 9'b111111111;
assign User[11][63] = 9'b111111111;
assign User[11][64] = 9'b111111111;
assign User[11][65] = 9'b111111111;
assign User[11][66] = 9'b111111111;
assign User[11][67] = 9'b111111111;
assign User[11][68] = 9'b111111111;
assign User[11][69] = 9'b111111111;
assign User[11][70] = 9'b111111111;
assign User[11][71] = 9'b111111111;
assign User[12][0] = 9'b111111111;
assign User[12][1] = 9'b111111111;
assign User[12][2] = 9'b111111111;
assign User[12][3] = 9'b111111111;
assign User[12][4] = 9'b111111111;
assign User[12][5] = 9'b111111111;
assign User[12][6] = 9'b111111111;
assign User[12][7] = 9'b111111111;
assign User[12][8] = 9'b111111111;
assign User[12][9] = 9'b111111111;
assign User[12][10] = 9'b111111111;
assign User[12][11] = 9'b111111111;
assign User[12][12] = 9'b111111111;
assign User[12][13] = 9'b111111111;
assign User[12][14] = 9'b111111111;
assign User[12][15] = 9'b111111111;
assign User[12][16] = 9'b111111111;
assign User[12][17] = 9'b111111111;
assign User[12][18] = 9'b111111111;
assign User[12][19] = 9'b111111111;
assign User[12][20] = 9'b111111111;
assign User[12][21] = 9'b111111111;
assign User[12][22] = 9'b111111111;
assign User[12][23] = 9'b111111111;
assign User[12][24] = 9'b111111111;
assign User[12][25] = 9'b111111111;
assign User[12][26] = 9'b111111111;
assign User[12][27] = 9'b111111111;
assign User[12][28] = 9'b111111111;
assign User[12][29] = 9'b111111111;
assign User[12][30] = 9'b111111111;
assign User[12][31] = 9'b111111111;
assign User[12][32] = 9'b111111111;
assign User[12][33] = 9'b111111111;
assign User[12][34] = 9'b111111111;
assign User[12][35] = 9'b111111111;
assign User[12][36] = 9'b111111111;
assign User[12][37] = 9'b111111111;
assign User[12][38] = 9'b111111111;
assign User[12][39] = 9'b111111111;
assign User[12][40] = 9'b111111111;
assign User[12][41] = 9'b111111111;
assign User[12][42] = 9'b111111111;
assign User[12][43] = 9'b111111111;
assign User[12][44] = 9'b111111111;
assign User[12][45] = 9'b111111111;
assign User[12][46] = 9'b111111111;
assign User[12][47] = 9'b111111111;
assign User[12][48] = 9'b111111111;
assign User[12][49] = 9'b111111111;
assign User[12][50] = 9'b111111111;
assign User[12][51] = 9'b111111111;
assign User[12][52] = 9'b111111111;
assign User[12][53] = 9'b111111111;
assign User[12][54] = 9'b111111111;
assign User[12][55] = 9'b111111111;
assign User[12][56] = 9'b111111111;
assign User[12][57] = 9'b111111111;
assign User[12][58] = 9'b111111111;
assign User[12][59] = 9'b111111111;
assign User[12][60] = 9'b111111111;
assign User[12][61] = 9'b111111111;
assign User[12][62] = 9'b111111111;
assign User[12][63] = 9'b111111111;
assign User[12][64] = 9'b111111111;
assign User[12][65] = 9'b111111111;
assign User[12][66] = 9'b111111111;
assign User[12][67] = 9'b111111111;
assign User[12][68] = 9'b111111111;
assign User[12][69] = 9'b111111111;
assign User[12][70] = 9'b111111111;
assign User[12][71] = 9'b111111111;
assign User[13][0] = 9'b111111111;
assign User[13][1] = 9'b111111111;
assign User[13][2] = 9'b111111111;
assign User[13][3] = 9'b111111111;
assign User[13][4] = 9'b111111111;
assign User[13][5] = 9'b111111111;
assign User[13][6] = 9'b111111111;
assign User[13][7] = 9'b111111111;
assign User[13][8] = 9'b111111111;
assign User[13][9] = 9'b111111111;
assign User[13][10] = 9'b111111111;
assign User[13][11] = 9'b111111111;
assign User[13][12] = 9'b111111111;
assign User[13][13] = 9'b111111111;
assign User[13][14] = 9'b111111111;
assign User[13][15] = 9'b111111111;
assign User[13][16] = 9'b111111111;
assign User[13][17] = 9'b111111111;
assign User[13][18] = 9'b111111111;
assign User[13][19] = 9'b111111111;
assign User[13][20] = 9'b111111111;
assign User[13][21] = 9'b111111111;
assign User[13][22] = 9'b111111111;
assign User[13][23] = 9'b111111111;
assign User[13][24] = 9'b111111111;
assign User[13][25] = 9'b111111111;
assign User[13][26] = 9'b111111111;
assign User[13][27] = 9'b111111111;
assign User[13][28] = 9'b111111111;
assign User[13][29] = 9'b111111111;
assign User[13][30] = 9'b111111111;
assign User[13][31] = 9'b111111111;
assign User[13][32] = 9'b111111111;
assign User[13][33] = 9'b111111111;
assign User[13][34] = 9'b111111111;
assign User[13][35] = 9'b111111111;
assign User[13][36] = 9'b111111111;
assign User[13][37] = 9'b111111111;
assign User[13][38] = 9'b111111111;
assign User[13][39] = 9'b111111111;
assign User[13][40] = 9'b111111111;
assign User[13][41] = 9'b111111111;
assign User[13][42] = 9'b111111111;
assign User[13][43] = 9'b111111111;
assign User[13][44] = 9'b111111111;
assign User[13][45] = 9'b111111111;
assign User[13][46] = 9'b111111111;
assign User[13][47] = 9'b111111111;
assign User[13][48] = 9'b111111111;
assign User[13][49] = 9'b111111111;
assign User[13][50] = 9'b111111111;
assign User[13][51] = 9'b111111111;
assign User[13][52] = 9'b111111111;
assign User[13][53] = 9'b111111111;
assign User[13][54] = 9'b111111111;
assign User[13][55] = 9'b111111111;
assign User[13][56] = 9'b111111111;
assign User[13][57] = 9'b111111111;
assign User[13][58] = 9'b111111111;
assign User[13][59] = 9'b111111111;
assign User[13][60] = 9'b111111111;
assign User[13][61] = 9'b111111111;
assign User[13][62] = 9'b111111111;
assign User[13][63] = 9'b111111111;
assign User[13][64] = 9'b111111111;
assign User[13][65] = 9'b111111111;
assign User[13][66] = 9'b111111111;
assign User[13][67] = 9'b111111111;
assign User[13][68] = 9'b111111111;
assign User[13][69] = 9'b111111111;
assign User[13][70] = 9'b111111111;
assign User[13][71] = 9'b111111111;
assign User[14][0] = 9'b111111111;
assign User[14][1] = 9'b111111111;
assign User[14][2] = 9'b111111111;
assign User[14][3] = 9'b111111111;
assign User[14][4] = 9'b111111111;
assign User[14][5] = 9'b111111111;
assign User[14][6] = 9'b111111111;
assign User[14][7] = 9'b111111111;
assign User[14][8] = 9'b111111111;
assign User[14][9] = 9'b111111111;
assign User[14][10] = 9'b111111111;
assign User[14][11] = 9'b111111111;
assign User[14][12] = 9'b111111111;
assign User[14][13] = 9'b111111111;
assign User[14][14] = 9'b111111111;
assign User[14][15] = 9'b111111111;
assign User[14][16] = 9'b111111111;
assign User[14][17] = 9'b111111111;
assign User[14][18] = 9'b111111111;
assign User[14][19] = 9'b111111111;
assign User[14][20] = 9'b111111111;
assign User[14][21] = 9'b111111111;
assign User[14][22] = 9'b111111111;
assign User[14][23] = 9'b111111111;
assign User[14][24] = 9'b111111111;
assign User[14][25] = 9'b111111111;
assign User[14][26] = 9'b111111111;
assign User[14][27] = 9'b111111111;
assign User[14][28] = 9'b111111111;
assign User[14][29] = 9'b111111111;
assign User[14][30] = 9'b111111111;
assign User[14][31] = 9'b111111111;
assign User[14][32] = 9'b111111111;
assign User[14][33] = 9'b111111111;
assign User[14][34] = 9'b111111111;
assign User[14][35] = 9'b111111111;
assign User[14][36] = 9'b111111111;
assign User[14][37] = 9'b111111111;
assign User[14][38] = 9'b111111111;
assign User[14][39] = 9'b111111111;
assign User[14][40] = 9'b111111111;
assign User[14][41] = 9'b111111111;
assign User[14][42] = 9'b101101101;
assign User[14][43] = 9'b111111111;
assign User[14][44] = 9'b111111111;
assign User[14][45] = 9'b111111111;
assign User[14][46] = 9'b111111111;
assign User[14][47] = 9'b111111111;
assign User[14][48] = 9'b111111111;
assign User[14][49] = 9'b111111111;
assign User[14][50] = 9'b111111111;
assign User[14][51] = 9'b111111111;
assign User[14][52] = 9'b111111111;
assign User[14][53] = 9'b111111111;
assign User[14][54] = 9'b111111111;
assign User[14][55] = 9'b111111111;
assign User[14][56] = 9'b111111111;
assign User[14][57] = 9'b111111111;
assign User[14][58] = 9'b111111111;
assign User[14][59] = 9'b111111111;
assign User[14][60] = 9'b111111111;
assign User[14][61] = 9'b111111111;
assign User[14][62] = 9'b111111111;
assign User[14][63] = 9'b111111111;
assign User[14][64] = 9'b111111111;
assign User[14][65] = 9'b111111111;
assign User[14][66] = 9'b111111111;
assign User[14][67] = 9'b111111111;
assign User[14][68] = 9'b111111111;
assign User[14][69] = 9'b111111111;
assign User[14][70] = 9'b111111111;
assign User[14][71] = 9'b111111111;
assign User[15][0] = 9'b111111111;
assign User[15][1] = 9'b111111111;
assign User[15][2] = 9'b111111111;
assign User[15][3] = 9'b111111111;
assign User[15][4] = 9'b111111111;
assign User[15][5] = 9'b111111111;
assign User[15][6] = 9'b111111111;
assign User[15][7] = 9'b111111111;
assign User[15][8] = 9'b111111111;
assign User[15][9] = 9'b111111111;
assign User[15][10] = 9'b111111111;
assign User[15][11] = 9'b111111111;
assign User[15][12] = 9'b111111111;
assign User[15][13] = 9'b111111111;
assign User[15][14] = 9'b111111111;
assign User[15][15] = 9'b111111111;
assign User[15][16] = 9'b111111111;
assign User[15][17] = 9'b111111111;
assign User[15][18] = 9'b111111111;
assign User[15][19] = 9'b111111111;
assign User[15][20] = 9'b111111111;
assign User[15][21] = 9'b111111111;
assign User[15][22] = 9'b111111111;
assign User[15][23] = 9'b111111111;
assign User[15][24] = 9'b111111111;
assign User[15][25] = 9'b111111111;
assign User[15][26] = 9'b101101101;
assign User[15][27] = 9'b100100100;
assign User[15][28] = 9'b100100100;
assign User[15][29] = 9'b110010010;
assign User[15][30] = 9'b111111111;
assign User[15][31] = 9'b101101101;
assign User[15][32] = 9'b100100100;
assign User[15][33] = 9'b100100100;
assign User[15][34] = 9'b110110110;
assign User[15][35] = 9'b111111111;
assign User[15][36] = 9'b101101101;
assign User[15][37] = 9'b100100100;
assign User[15][38] = 9'b111111111;
assign User[15][39] = 9'b111111111;
assign User[15][40] = 9'b111111111;
assign User[15][41] = 9'b101101101;
assign User[15][42] = 9'b100100100;
assign User[15][43] = 9'b101101101;
assign User[15][44] = 9'b111111111;
assign User[15][45] = 9'b111111111;
assign User[15][46] = 9'b111111111;
assign User[15][47] = 9'b111111111;
assign User[15][48] = 9'b110110110;
assign User[15][49] = 9'b100100100;
assign User[15][50] = 9'b100100100;
assign User[15][51] = 9'b110010001;
assign User[15][52] = 9'b111111111;
assign User[15][53] = 9'b101101101;
assign User[15][54] = 9'b100100100;
assign User[15][55] = 9'b100100100;
assign User[15][56] = 9'b110010010;
assign User[15][57] = 9'b111111111;
assign User[15][58] = 9'b110010001;
assign User[15][59] = 9'b101101101;
assign User[15][60] = 9'b111111111;
assign User[15][61] = 9'b111111111;
assign User[15][62] = 9'b111111111;
assign User[15][63] = 9'b101001001;
assign User[15][64] = 9'b100100100;
assign User[15][65] = 9'b101101101;
assign User[15][66] = 9'b111111111;
assign User[15][67] = 9'b111111111;
assign User[15][68] = 9'b111111111;
assign User[15][69] = 9'b111111111;
assign User[15][70] = 9'b111111111;
assign User[15][71] = 9'b111111111;
assign User[16][0] = 9'b111111111;
assign User[16][1] = 9'b111111111;
assign User[16][2] = 9'b111111111;
assign User[16][3] = 9'b111111111;
assign User[16][4] = 9'b111111111;
assign User[16][5] = 9'b111111111;
assign User[16][6] = 9'b111111111;
assign User[16][7] = 9'b111111111;
assign User[16][8] = 9'b111111111;
assign User[16][9] = 9'b111111111;
assign User[16][10] = 9'b111111111;
assign User[16][11] = 9'b111111111;
assign User[16][12] = 9'b111111111;
assign User[16][13] = 9'b111111111;
assign User[16][14] = 9'b111111111;
assign User[16][15] = 9'b111111111;
assign User[16][16] = 9'b111111111;
assign User[16][17] = 9'b111111111;
assign User[16][18] = 9'b111111111;
assign User[16][19] = 9'b111111111;
assign User[16][20] = 9'b111111111;
assign User[16][21] = 9'b111111111;
assign User[16][22] = 9'b111111111;
assign User[16][23] = 9'b111111111;
assign User[16][24] = 9'b111111111;
assign User[16][25] = 9'b111111111;
assign User[16][26] = 9'b101001000;
assign User[16][27] = 9'b110010010;
assign User[16][28] = 9'b101101101;
assign User[16][29] = 9'b100100100;
assign User[16][30] = 9'b111111111;
assign User[16][31] = 9'b100100100;
assign User[16][32] = 9'b110110110;
assign User[16][33] = 9'b110010001;
assign User[16][34] = 9'b101001001;
assign User[16][35] = 9'b111111111;
assign User[16][36] = 9'b101101101;
assign User[16][37] = 9'b100100100;
assign User[16][38] = 9'b111111111;
assign User[16][39] = 9'b111111111;
assign User[16][40] = 9'b110010010;
assign User[16][41] = 9'b101001001;
assign User[16][42] = 9'b110110110;
assign User[16][43] = 9'b101101101;
assign User[16][44] = 9'b111111111;
assign User[16][45] = 9'b111111111;
assign User[16][46] = 9'b111111111;
assign User[16][47] = 9'b111111111;
assign User[16][48] = 9'b101001000;
assign User[16][49] = 9'b101101101;
assign User[16][50] = 9'b101001001;
assign User[16][51] = 9'b110010001;
assign User[16][52] = 9'b111111111;
assign User[16][53] = 9'b101001000;
assign User[16][54] = 9'b110010010;
assign User[16][55] = 9'b101101101;
assign User[16][56] = 9'b100100100;
assign User[16][57] = 9'b111111111;
assign User[16][58] = 9'b101101101;
assign User[16][59] = 9'b101101101;
assign User[16][60] = 9'b111111111;
assign User[16][61] = 9'b111111111;
assign User[16][62] = 9'b101101101;
assign User[16][63] = 9'b101101101;
assign User[16][64] = 9'b111111111;
assign User[16][65] = 9'b100100100;
assign User[16][66] = 9'b111111111;
assign User[16][67] = 9'b111111111;
assign User[16][68] = 9'b111111111;
assign User[16][69] = 9'b111111111;
assign User[16][70] = 9'b111111111;
assign User[16][71] = 9'b111111111;
assign User[17][0] = 9'b111111111;
assign User[17][1] = 9'b111111111;
assign User[17][2] = 9'b111111111;
assign User[17][3] = 9'b111111111;
assign User[17][4] = 9'b111111111;
assign User[17][5] = 9'b111111111;
assign User[17][6] = 9'b111111111;
assign User[17][7] = 9'b111111111;
assign User[17][8] = 9'b111111111;
assign User[17][9] = 9'b111111111;
assign User[17][10] = 9'b111111111;
assign User[17][11] = 9'b111111111;
assign User[17][12] = 9'b111111111;
assign User[17][13] = 9'b111111111;
assign User[17][14] = 9'b111111111;
assign User[17][15] = 9'b111111111;
assign User[17][16] = 9'b111111111;
assign User[17][17] = 9'b111111111;
assign User[17][18] = 9'b111111111;
assign User[17][19] = 9'b111111111;
assign User[17][20] = 9'b111111111;
assign User[17][21] = 9'b111111111;
assign User[17][22] = 9'b111111111;
assign User[17][23] = 9'b111111111;
assign User[17][24] = 9'b111111111;
assign User[17][25] = 9'b111111111;
assign User[17][26] = 9'b101101101;
assign User[17][27] = 9'b100100100;
assign User[17][28] = 9'b101001001;
assign User[17][29] = 9'b110010001;
assign User[17][30] = 9'b110010010;
assign User[17][31] = 9'b101001000;
assign User[17][32] = 9'b111111111;
assign User[17][33] = 9'b111111111;
assign User[17][34] = 9'b100100100;
assign User[17][35] = 9'b111111111;
assign User[17][36] = 9'b111111111;
assign User[17][37] = 9'b100100100;
assign User[17][38] = 9'b111111111;
assign User[17][39] = 9'b111111111;
assign User[17][40] = 9'b111111111;
assign User[17][41] = 9'b101001001;
assign User[17][42] = 9'b100100100;
assign User[17][43] = 9'b101001001;
assign User[17][44] = 9'b111111111;
assign User[17][45] = 9'b101101101;
assign User[17][46] = 9'b101101101;
assign User[17][47] = 9'b110010001;
assign User[17][48] = 9'b100100100;
assign User[17][49] = 9'b101101101;
assign User[17][50] = 9'b101001000;
assign User[17][51] = 9'b110010001;
assign User[17][52] = 9'b111111111;
assign User[17][53] = 9'b101101101;
assign User[17][54] = 9'b100100100;
assign User[17][55] = 9'b101001001;
assign User[17][56] = 9'b110010001;
assign User[17][57] = 9'b111111111;
assign User[17][58] = 9'b111111111;
assign User[17][59] = 9'b101101101;
assign User[17][60] = 9'b101101101;
assign User[17][61] = 9'b111111111;
assign User[17][62] = 9'b101101101;
assign User[17][63] = 9'b101101101;
assign User[17][64] = 9'b111111111;
assign User[17][65] = 9'b100100100;
assign User[17][66] = 9'b110010010;
assign User[17][67] = 9'b111111111;
assign User[17][68] = 9'b111111111;
assign User[17][69] = 9'b111111111;
assign User[17][70] = 9'b111111111;
assign User[17][71] = 9'b111111111;
assign User[18][0] = 9'b111111111;
assign User[18][1] = 9'b111111111;
assign User[18][2] = 9'b111111111;
assign User[18][3] = 9'b111111111;
assign User[18][4] = 9'b111111111;
assign User[18][5] = 9'b111111111;
assign User[18][6] = 9'b111111111;
assign User[18][7] = 9'b111111111;
assign User[18][8] = 9'b111111111;
assign User[18][9] = 9'b111111111;
assign User[18][10] = 9'b111111111;
assign User[18][11] = 9'b111111111;
assign User[18][12] = 9'b111111111;
assign User[18][13] = 9'b111111111;
assign User[18][14] = 9'b111111111;
assign User[18][15] = 9'b111111111;
assign User[18][16] = 9'b111111111;
assign User[18][17] = 9'b111111111;
assign User[18][18] = 9'b111111111;
assign User[18][19] = 9'b111111111;
assign User[18][20] = 9'b111111111;
assign User[18][21] = 9'b111111111;
assign User[18][22] = 9'b111111111;
assign User[18][23] = 9'b111111111;
assign User[18][24] = 9'b111111111;
assign User[18][25] = 9'b111111111;
assign User[18][26] = 9'b111111111;
assign User[18][27] = 9'b101101101;
assign User[18][28] = 9'b110010001;
assign User[18][29] = 9'b111111111;
assign User[18][30] = 9'b110110110;
assign User[18][31] = 9'b101001000;
assign User[18][32] = 9'b111111111;
assign User[18][33] = 9'b111111111;
assign User[18][34] = 9'b100100100;
assign User[18][35] = 9'b111111111;
assign User[18][36] = 9'b111111111;
assign User[18][37] = 9'b100100100;
assign User[18][38] = 9'b111111111;
assign User[18][39] = 9'b111111111;
assign User[18][40] = 9'b101101101;
assign User[18][41] = 9'b110010001;
assign User[18][42] = 9'b111111111;
assign User[18][43] = 9'b101101101;
assign User[18][44] = 9'b101101101;
assign User[18][45] = 9'b110010001;
assign User[18][46] = 9'b101001001;
assign User[18][47] = 9'b101101101;
assign User[18][48] = 9'b100100100;
assign User[18][49] = 9'b110110110;
assign User[18][50] = 9'b110010001;
assign User[18][51] = 9'b101001000;
assign User[18][52] = 9'b111111111;
assign User[18][53] = 9'b111111111;
assign User[18][54] = 9'b101101101;
assign User[18][55] = 9'b110010001;
assign User[18][56] = 9'b111111111;
assign User[18][57] = 9'b101101101;
assign User[18][58] = 9'b101001001;
assign User[18][59] = 9'b101001000;
assign User[18][60] = 9'b101001000;
assign User[18][61] = 9'b111111111;
assign User[18][62] = 9'b111111111;
assign User[18][63] = 9'b100100100;
assign User[18][64] = 9'b100100100;
assign User[18][65] = 9'b100100100;
assign User[18][66] = 9'b110110110;
assign User[18][67] = 9'b111111111;
assign User[18][68] = 9'b111111111;
assign User[18][69] = 9'b111111111;
assign User[18][70] = 9'b111111111;
assign User[18][71] = 9'b111111111;
assign User[19][0] = 9'b111111111;
assign User[19][1] = 9'b111111111;
assign User[19][2] = 9'b111111111;
assign User[19][3] = 9'b111111111;
assign User[19][4] = 9'b111111111;
assign User[19][5] = 9'b111111111;
assign User[19][6] = 9'b111111111;
assign User[19][7] = 9'b111111111;
assign User[19][8] = 9'b111111111;
assign User[19][9] = 9'b111111111;
assign User[19][10] = 9'b111111111;
assign User[19][11] = 9'b111111111;
assign User[19][12] = 9'b111111111;
assign User[19][13] = 9'b111111111;
assign User[19][14] = 9'b111111111;
assign User[19][15] = 9'b111111111;
assign User[19][16] = 9'b111111111;
assign User[19][17] = 9'b111111111;
assign User[19][18] = 9'b111111111;
assign User[19][19] = 9'b111111111;
assign User[19][20] = 9'b111111111;
assign User[19][21] = 9'b111111111;
assign User[19][22] = 9'b111111111;
assign User[19][23] = 9'b111111111;
assign User[19][24] = 9'b111111111;
assign User[19][25] = 9'b111111111;
assign User[19][26] = 9'b100100100;
assign User[19][27] = 9'b100100100;
assign User[19][28] = 9'b101101101;
assign User[19][29] = 9'b101001001;
assign User[19][30] = 9'b111111111;
assign User[19][31] = 9'b101001001;
assign User[19][32] = 9'b110010001;
assign User[19][33] = 9'b101101101;
assign User[19][34] = 9'b101101101;
assign User[19][35] = 9'b111111111;
assign User[19][36] = 9'b110110110;
assign User[19][37] = 9'b100000000;
assign User[19][38] = 9'b111111111;
assign User[19][39] = 9'b111111111;
assign User[19][40] = 9'b101101101;
assign User[19][41] = 9'b101101101;
assign User[19][42] = 9'b111111111;
assign User[19][43] = 9'b101101101;
assign User[19][44] = 9'b110010001;
assign User[19][45] = 9'b111111111;
assign User[19][46] = 9'b111111111;
assign User[19][47] = 9'b111111111;
assign User[19][48] = 9'b101001001;
assign User[19][49] = 9'b110010001;
assign User[19][50] = 9'b101101101;
assign User[19][51] = 9'b101101101;
assign User[19][52] = 9'b111111111;
assign User[19][53] = 9'b100100100;
assign User[19][54] = 9'b100100100;
assign User[19][55] = 9'b101101101;
assign User[19][56] = 9'b101001000;
assign User[19][57] = 9'b111111111;
assign User[19][58] = 9'b111111111;
assign User[19][59] = 9'b100100100;
assign User[19][60] = 9'b100100100;
assign User[19][61] = 9'b110110110;
assign User[19][62] = 9'b111111111;
assign User[19][63] = 9'b111111111;
assign User[19][64] = 9'b110010010;
assign User[19][65] = 9'b101001001;
assign User[19][66] = 9'b111111111;
assign User[19][67] = 9'b111111111;
assign User[19][68] = 9'b111111111;
assign User[19][69] = 9'b111111111;
assign User[19][70] = 9'b111111111;
assign User[19][71] = 9'b111111111;
assign User[20][0] = 9'b111111111;
assign User[20][1] = 9'b111111111;
assign User[20][2] = 9'b111111111;
assign User[20][3] = 9'b111111111;
assign User[20][4] = 9'b111111111;
assign User[20][5] = 9'b111111111;
assign User[20][6] = 9'b111111111;
assign User[20][7] = 9'b111111111;
assign User[20][8] = 9'b111111111;
assign User[20][9] = 9'b111111111;
assign User[20][10] = 9'b111111111;
assign User[20][11] = 9'b111111111;
assign User[20][12] = 9'b111111111;
assign User[20][13] = 9'b111111111;
assign User[20][14] = 9'b111111111;
assign User[20][15] = 9'b111111111;
assign User[20][16] = 9'b111111111;
assign User[20][17] = 9'b111111111;
assign User[20][18] = 9'b111111111;
assign User[20][19] = 9'b111111111;
assign User[20][20] = 9'b111111111;
assign User[20][21] = 9'b111111111;
assign User[20][22] = 9'b111111111;
assign User[20][23] = 9'b111111111;
assign User[20][24] = 9'b111111111;
assign User[20][25] = 9'b111111111;
assign User[20][26] = 9'b110010001;
assign User[20][27] = 9'b101101101;
assign User[20][28] = 9'b101101101;
assign User[20][29] = 9'b101101101;
assign User[20][30] = 9'b111111111;
assign User[20][31] = 9'b111111111;
assign User[20][32] = 9'b101101101;
assign User[20][33] = 9'b110010001;
assign User[20][34] = 9'b111111111;
assign User[20][35] = 9'b111111111;
assign User[20][36] = 9'b110110110;
assign User[20][37] = 9'b101101101;
assign User[20][38] = 9'b110110110;
assign User[20][39] = 9'b111111111;
assign User[20][40] = 9'b111111111;
assign User[20][41] = 9'b101101101;
assign User[20][42] = 9'b101101101;
assign User[20][43] = 9'b110010010;
assign User[20][44] = 9'b111111111;
assign User[20][45] = 9'b111111111;
assign User[20][46] = 9'b111111111;
assign User[20][47] = 9'b111111111;
assign User[20][48] = 9'b111111111;
assign User[20][49] = 9'b101101101;
assign User[20][50] = 9'b110010001;
assign User[20][51] = 9'b111111111;
assign User[20][52] = 9'b111111111;
assign User[20][53] = 9'b110010001;
assign User[20][54] = 9'b101101101;
assign User[20][55] = 9'b101101101;
assign User[20][56] = 9'b101101101;
assign User[20][57] = 9'b111111111;
assign User[20][58] = 9'b111111111;
assign User[20][59] = 9'b101101101;
assign User[20][60] = 9'b101101101;
assign User[20][61] = 9'b111111111;
assign User[20][62] = 9'b111111111;
assign User[20][63] = 9'b101101101;
assign User[20][64] = 9'b101001001;
assign User[20][65] = 9'b110110110;
assign User[20][66] = 9'b111111111;
assign User[20][67] = 9'b111111111;
assign User[20][68] = 9'b111111111;
assign User[20][69] = 9'b111111111;
assign User[20][70] = 9'b111111111;
assign User[20][71] = 9'b111111111;
assign User[21][0] = 9'b111111111;
assign User[21][1] = 9'b111111111;
assign User[21][2] = 9'b111111111;
assign User[21][3] = 9'b111111111;
assign User[21][4] = 9'b111111111;
assign User[21][5] = 9'b111111111;
assign User[21][6] = 9'b111111111;
assign User[21][7] = 9'b111111111;
assign User[21][8] = 9'b111111111;
assign User[21][9] = 9'b111111111;
assign User[21][10] = 9'b111111111;
assign User[21][11] = 9'b111111111;
assign User[21][12] = 9'b111111111;
assign User[21][13] = 9'b111111111;
assign User[21][14] = 9'b111111111;
assign User[21][15] = 9'b111111111;
assign User[21][16] = 9'b111111111;
assign User[21][17] = 9'b111111111;
assign User[21][18] = 9'b111111111;
assign User[21][19] = 9'b111111111;
assign User[21][20] = 9'b111111111;
assign User[21][21] = 9'b111111111;
assign User[21][22] = 9'b111111111;
assign User[21][23] = 9'b111111111;
assign User[21][24] = 9'b111111111;
assign User[21][25] = 9'b111111111;
assign User[21][26] = 9'b111111111;
assign User[21][27] = 9'b111111111;
assign User[21][28] = 9'b111111111;
assign User[21][29] = 9'b111111111;
assign User[21][30] = 9'b111111111;
assign User[21][31] = 9'b111111111;
assign User[21][32] = 9'b111111111;
assign User[21][33] = 9'b111111111;
assign User[21][34] = 9'b111111111;
assign User[21][35] = 9'b111111111;
assign User[21][36] = 9'b111111111;
assign User[21][37] = 9'b111111111;
assign User[21][38] = 9'b111111111;
assign User[21][39] = 9'b111111111;
assign User[21][40] = 9'b111111111;
assign User[21][41] = 9'b111111111;
assign User[21][42] = 9'b111111111;
assign User[21][43] = 9'b111111111;
assign User[21][44] = 9'b111111111;
assign User[21][45] = 9'b111111111;
assign User[21][46] = 9'b111111111;
assign User[21][47] = 9'b111111111;
assign User[21][48] = 9'b111111111;
assign User[21][49] = 9'b111111111;
assign User[21][50] = 9'b111111111;
assign User[21][51] = 9'b111111111;
assign User[21][52] = 9'b111111111;
assign User[21][53] = 9'b111111111;
assign User[21][54] = 9'b111111111;
assign User[21][55] = 9'b111111111;
assign User[21][56] = 9'b111111111;
assign User[21][57] = 9'b111111111;
assign User[21][58] = 9'b111111111;
assign User[21][59] = 9'b111111111;
assign User[21][60] = 9'b111111111;
assign User[21][61] = 9'b111111111;
assign User[21][62] = 9'b111111111;
assign User[21][63] = 9'b101101101;
assign User[21][64] = 9'b110110110;
assign User[21][65] = 9'b111111111;
assign User[21][66] = 9'b111111111;
assign User[21][67] = 9'b111111111;
assign User[21][68] = 9'b111111111;
assign User[21][69] = 9'b111111111;
assign User[21][70] = 9'b111111111;
assign User[21][71] = 9'b111111111;
assign User[22][0] = 9'b111111111;
assign User[22][1] = 9'b111111111;
assign User[22][2] = 9'b111111111;
assign User[22][3] = 9'b111111111;
assign User[22][4] = 9'b111111111;
assign User[22][5] = 9'b111111111;
assign User[22][6] = 9'b111111111;
assign User[22][7] = 9'b111111111;
assign User[22][8] = 9'b111111111;
assign User[22][9] = 9'b111111111;
assign User[22][10] = 9'b111111111;
assign User[22][11] = 9'b111111111;
assign User[22][12] = 9'b111111111;
assign User[22][13] = 9'b111111111;
assign User[22][14] = 9'b111111111;
assign User[22][15] = 9'b111111111;
assign User[22][16] = 9'b111111111;
assign User[22][17] = 9'b111111111;
assign User[22][18] = 9'b111111111;
assign User[22][19] = 9'b111111111;
assign User[22][20] = 9'b111111111;
assign User[22][21] = 9'b111111111;
assign User[22][22] = 9'b111111111;
assign User[22][23] = 9'b111111111;
assign User[22][24] = 9'b111111111;
assign User[22][25] = 9'b111111111;
assign User[22][26] = 9'b111111111;
assign User[22][27] = 9'b111111111;
assign User[22][28] = 9'b111111111;
assign User[22][29] = 9'b111111111;
assign User[22][30] = 9'b111111111;
assign User[22][31] = 9'b111111111;
assign User[22][32] = 9'b111111111;
assign User[22][33] = 9'b111111111;
assign User[22][34] = 9'b111111111;
assign User[22][35] = 9'b111111111;
assign User[22][36] = 9'b111111111;
assign User[22][37] = 9'b111111111;
assign User[22][38] = 9'b111111111;
assign User[22][39] = 9'b111111111;
assign User[22][40] = 9'b111111111;
assign User[22][41] = 9'b111111111;
assign User[22][42] = 9'b111111111;
assign User[22][43] = 9'b111111111;
assign User[22][44] = 9'b111111111;
assign User[22][45] = 9'b111111111;
assign User[22][46] = 9'b111111111;
assign User[22][47] = 9'b111111111;
assign User[22][48] = 9'b111111111;
assign User[22][49] = 9'b111111111;
assign User[22][50] = 9'b111111111;
assign User[22][51] = 9'b111111111;
assign User[22][52] = 9'b111111111;
assign User[22][53] = 9'b111111111;
assign User[22][54] = 9'b111111111;
assign User[22][55] = 9'b111111111;
assign User[22][56] = 9'b111111111;
assign User[22][57] = 9'b111111111;
assign User[22][58] = 9'b111111111;
assign User[22][59] = 9'b111111111;
assign User[22][60] = 9'b111111111;
assign User[22][61] = 9'b111111111;
assign User[22][62] = 9'b111111111;
assign User[22][63] = 9'b111111111;
assign User[22][64] = 9'b111111111;
assign User[22][65] = 9'b111111111;
assign User[22][66] = 9'b111111111;
assign User[22][67] = 9'b111111111;
assign User[22][68] = 9'b111111111;
assign User[22][69] = 9'b111111111;
assign User[22][70] = 9'b111111111;
assign User[22][71] = 9'b111111111;
assign User[23][0] = 9'b111111111;
assign User[23][1] = 9'b111111111;
assign User[23][2] = 9'b111111111;
assign User[23][3] = 9'b111111111;
assign User[23][4] = 9'b111111111;
assign User[23][5] = 9'b111111111;
assign User[23][6] = 9'b111111111;
assign User[23][7] = 9'b111111111;
assign User[23][8] = 9'b111111111;
assign User[23][9] = 9'b111111111;
assign User[23][10] = 9'b111111111;
assign User[23][11] = 9'b111111111;
assign User[23][12] = 9'b111111111;
assign User[23][13] = 9'b111111111;
assign User[23][14] = 9'b111111111;
assign User[23][15] = 9'b111111111;
assign User[23][16] = 9'b111111111;
assign User[23][17] = 9'b111111111;
assign User[23][18] = 9'b111111111;
assign User[23][19] = 9'b111111111;
assign User[23][20] = 9'b111111111;
assign User[23][21] = 9'b111111111;
assign User[23][22] = 9'b111111111;
assign User[23][23] = 9'b111111111;
assign User[23][24] = 9'b111111111;
assign User[23][25] = 9'b111111111;
assign User[23][26] = 9'b111111111;
assign User[23][27] = 9'b111111111;
assign User[23][28] = 9'b111111111;
assign User[23][29] = 9'b111111111;
assign User[23][30] = 9'b111111111;
assign User[23][31] = 9'b111111111;
assign User[23][32] = 9'b111111111;
assign User[23][33] = 9'b111111111;
assign User[23][34] = 9'b111111111;
assign User[23][35] = 9'b111111111;
assign User[23][36] = 9'b111111111;
assign User[23][37] = 9'b111111111;
assign User[23][38] = 9'b111111111;
assign User[23][39] = 9'b111111111;
assign User[23][40] = 9'b111111111;
assign User[23][41] = 9'b111111111;
assign User[23][42] = 9'b111111111;
assign User[23][43] = 9'b111111111;
assign User[23][44] = 9'b111111111;
assign User[23][45] = 9'b111111111;
assign User[23][46] = 9'b111111111;
assign User[23][47] = 9'b111111111;
assign User[23][48] = 9'b111111111;
assign User[23][49] = 9'b111111111;
assign User[23][50] = 9'b111111111;
assign User[23][51] = 9'b111111111;
assign User[23][52] = 9'b111111111;
assign User[23][53] = 9'b111111111;
assign User[23][54] = 9'b111111111;
assign User[23][55] = 9'b111111111;
assign User[23][56] = 9'b111111111;
assign User[23][57] = 9'b111111111;
assign User[23][58] = 9'b111111111;
assign User[23][59] = 9'b111111111;
assign User[23][60] = 9'b111111111;
assign User[23][61] = 9'b111111111;
assign User[23][62] = 9'b111111111;
assign User[23][63] = 9'b111111111;
assign User[23][64] = 9'b111111111;
assign User[23][65] = 9'b111111111;
assign User[23][66] = 9'b111111111;
assign User[23][67] = 9'b111111111;
assign User[23][68] = 9'b111111111;
assign User[23][69] = 9'b111111111;
assign User[23][70] = 9'b111111111;
assign User[23][71] = 9'b111111111;
assign User[24][0] = 9'b111111111;
assign User[24][1] = 9'b111111111;
assign User[24][2] = 9'b111111111;
assign User[24][3] = 9'b111111111;
assign User[24][4] = 9'b111111111;
assign User[24][5] = 9'b111111111;
assign User[24][6] = 9'b111111111;
assign User[24][7] = 9'b111111111;
assign User[24][8] = 9'b111111111;
assign User[24][9] = 9'b111111111;
assign User[24][10] = 9'b111111111;
assign User[24][11] = 9'b111111111;
assign User[24][12] = 9'b111111111;
assign User[24][13] = 9'b111111111;
assign User[24][14] = 9'b111111111;
assign User[24][15] = 9'b111111111;
assign User[24][16] = 9'b111111111;
assign User[24][17] = 9'b111111111;
assign User[24][18] = 9'b111111111;
assign User[24][19] = 9'b111111111;
assign User[24][20] = 9'b111111111;
assign User[24][21] = 9'b111111111;
assign User[24][22] = 9'b111111111;
assign User[24][23] = 9'b111111111;
assign User[24][24] = 9'b111111111;
assign User[24][25] = 9'b111111111;
assign User[24][26] = 9'b111111111;
assign User[24][27] = 9'b111111111;
assign User[24][28] = 9'b111111111;
assign User[24][29] = 9'b111111111;
assign User[24][30] = 9'b111111111;
assign User[24][31] = 9'b111111111;
assign User[24][32] = 9'b111111111;
assign User[24][33] = 9'b111111111;
assign User[24][34] = 9'b111111111;
assign User[24][35] = 9'b111111111;
assign User[24][36] = 9'b111111111;
assign User[24][37] = 9'b111111111;
assign User[24][38] = 9'b111111111;
assign User[24][39] = 9'b111111111;
assign User[24][40] = 9'b111111111;
assign User[24][41] = 9'b111111111;
assign User[24][42] = 9'b111111111;
assign User[24][43] = 9'b111111111;
assign User[24][44] = 9'b111111111;
assign User[24][45] = 9'b111111111;
assign User[24][46] = 9'b111111111;
assign User[24][47] = 9'b111111111;
assign User[24][48] = 9'b111111111;
assign User[24][49] = 9'b111111111;
assign User[24][50] = 9'b111111111;
assign User[24][51] = 9'b111111111;
assign User[24][52] = 9'b111111111;
assign User[24][53] = 9'b111111111;
assign User[24][54] = 9'b111111111;
assign User[24][55] = 9'b111111111;
assign User[24][56] = 9'b111111111;
assign User[24][57] = 9'b111111111;
assign User[24][58] = 9'b111111111;
assign User[24][59] = 9'b111111111;
assign User[24][60] = 9'b111111111;
assign User[24][61] = 9'b111111111;
assign User[24][62] = 9'b111111111;
assign User[24][63] = 9'b111111111;
assign User[24][64] = 9'b111111111;
assign User[24][65] = 9'b111111111;
assign User[24][66] = 9'b111111111;
assign User[24][67] = 9'b111111111;
assign User[24][68] = 9'b111111111;
assign User[24][69] = 9'b111111111;
assign User[24][70] = 9'b111111111;
assign User[24][71] = 9'b111111111;
//Total de Lineas = 1800

endmodule
