`timescale 1ns / 1ps
module Boton_Exit (
input enable,
input clock,
input [9:0] posx, posy,
input [9:0] hcount,
input [9:0] vcount,
output reg[2:0] red,
output reg[2:0] green,
output reg[1:0] blue,
output reg data);

always @(posedge clock)
begin
	if(enable)
	begin
		if(hcount >= posx & hcount < posx + RESOLUCION_X & vcount >= posy & vcount < posy + RESOLUCION_Y)
		begin
			if (Boton[vcount - posy][hcount - posx][8] == 1'b1)
			begin
				red   <= Boton[vcount- posy][hcount- posx][7:5];
				green <= Boton[vcount- posy][hcount- posx][4:2];
            blue 	<= Boton[vcount- posy][hcount- posx][1:0];
				data  <= 1'b1;
			end
			else
				data <= 0;
			end
		else
		data <= 0;
	end
	end
parameter RESOLUCION_X = 50;
parameter RESOLUCION_Y = 50;
wire [9:0] Boton[RESOLUCION_Y - 1'b1 : 0][RESOLUCION_X - 1'b1 : 0];
assign Boton[1][20] = 9'b101001001;
assign Boton[1][21] = 9'b101000100;
assign Boton[1][22] = 9'b100100100;
assign Boton[1][23] = 9'b100100000;
assign Boton[1][24] = 9'b100100100;
assign Boton[1][25] = 9'b100100100;
assign Boton[1][26] = 9'b100100100;
assign Boton[1][27] = 9'b100100100;
assign Boton[1][28] = 9'b101001001;
assign Boton[2][17] = 9'b100100100;
assign Boton[2][18] = 9'b100100100;
assign Boton[2][19] = 9'b100100100;
assign Boton[2][20] = 9'b100100100;
assign Boton[2][21] = 9'b100100100;
assign Boton[2][22] = 9'b100000000;
assign Boton[2][23] = 9'b100000000;
assign Boton[2][24] = 9'b100000100;
assign Boton[2][25] = 9'b100000100;
assign Boton[2][26] = 9'b100000000;
assign Boton[2][27] = 9'b100000000;
assign Boton[2][28] = 9'b100100100;
assign Boton[2][29] = 9'b100100100;
assign Boton[2][30] = 9'b100100100;
assign Boton[2][31] = 9'b100100100;
assign Boton[3][15] = 9'b100100100;
assign Boton[3][16] = 9'b100100100;
assign Boton[3][17] = 9'b100000000;
assign Boton[3][18] = 9'b100000000;
assign Boton[3][19] = 9'b100000100;
assign Boton[3][20] = 9'b100000100;
assign Boton[3][21] = 9'b100001001;
assign Boton[3][22] = 9'b100001001;
assign Boton[3][23] = 9'b100001001;
assign Boton[3][24] = 9'b100001001;
assign Boton[3][25] = 9'b100001001;
assign Boton[3][26] = 9'b100001001;
assign Boton[3][27] = 9'b100000101;
assign Boton[3][28] = 9'b100000100;
assign Boton[3][29] = 9'b100000100;
assign Boton[3][30] = 9'b100000000;
assign Boton[3][31] = 9'b100100000;
assign Boton[3][32] = 9'b100100000;
assign Boton[3][33] = 9'b100100100;
assign Boton[3][34] = 9'b101001000;
assign Boton[4][13] = 9'b100100100;
assign Boton[4][14] = 9'b100100100;
assign Boton[4][15] = 9'b100100000;
assign Boton[4][16] = 9'b100000100;
assign Boton[4][17] = 9'b100001001;
assign Boton[4][18] = 9'b100001001;
assign Boton[4][19] = 9'b100001001;
assign Boton[4][20] = 9'b100101001;
assign Boton[4][21] = 9'b100101001;
assign Boton[4][22] = 9'b100001001;
assign Boton[4][23] = 9'b100001001;
assign Boton[4][24] = 9'b100001001;
assign Boton[4][25] = 9'b100001001;
assign Boton[4][26] = 9'b100001001;
assign Boton[4][27] = 9'b100001001;
assign Boton[4][28] = 9'b100001001;
assign Boton[4][29] = 9'b100001001;
assign Boton[4][30] = 9'b100001001;
assign Boton[4][31] = 9'b100000101;
assign Boton[4][32] = 9'b100000100;
assign Boton[4][33] = 9'b100000000;
assign Boton[4][34] = 9'b100100000;
assign Boton[4][35] = 9'b100100100;
assign Boton[4][36] = 9'b101001101;
assign Boton[5][12] = 9'b100100100;
assign Boton[5][13] = 9'b100100000;
assign Boton[5][14] = 9'b100000100;
assign Boton[5][15] = 9'b100001001;
assign Boton[5][16] = 9'b100001001;
assign Boton[5][17] = 9'b100001001;
assign Boton[5][18] = 9'b100000101;
assign Boton[5][19] = 9'b100001001;
assign Boton[5][20] = 9'b100001101;
assign Boton[5][21] = 9'b100001110;
assign Boton[5][22] = 9'b100010010;
assign Boton[5][23] = 9'b100010010;
assign Boton[5][24] = 9'b100010010;
assign Boton[5][25] = 9'b100010010;
assign Boton[5][26] = 9'b100010010;
assign Boton[5][27] = 9'b100010010;
assign Boton[5][28] = 9'b100010010;
assign Boton[5][29] = 9'b100001001;
assign Boton[5][30] = 9'b100001001;
assign Boton[5][31] = 9'b100001101;
assign Boton[5][32] = 9'b100001001;
assign Boton[5][33] = 9'b100001001;
assign Boton[5][34] = 9'b100000100;
assign Boton[5][35] = 9'b100000000;
assign Boton[5][36] = 9'b100100100;
assign Boton[5][37] = 9'b101001001;
assign Boton[6][10] = 9'b100100100;
assign Boton[6][11] = 9'b100100100;
assign Boton[6][12] = 9'b100000000;
assign Boton[6][13] = 9'b100000100;
assign Boton[6][14] = 9'b100001001;
assign Boton[6][15] = 9'b100101001;
assign Boton[6][16] = 9'b100101001;
assign Boton[6][17] = 9'b100001101;
assign Boton[6][18] = 9'b100001001;
assign Boton[6][19] = 9'b100001001;
assign Boton[6][20] = 9'b100010011;
assign Boton[6][21] = 9'b100010010;
assign Boton[6][22] = 9'b100001101;
assign Boton[6][23] = 9'b100001001;
assign Boton[6][24] = 9'b100001001;
assign Boton[6][25] = 9'b100001001;
assign Boton[6][26] = 9'b100001001;
assign Boton[6][27] = 9'b100001001;
assign Boton[6][28] = 9'b100001001;
assign Boton[6][29] = 9'b100000100;
assign Boton[6][30] = 9'b100000101;
assign Boton[6][31] = 9'b100001101;
assign Boton[6][32] = 9'b100001101;
assign Boton[6][33] = 9'b100001101;
assign Boton[6][34] = 9'b100001001;
assign Boton[6][35] = 9'b100000100;
assign Boton[6][36] = 9'b100000000;
assign Boton[6][37] = 9'b100100100;
assign Boton[6][38] = 9'b100100100;
assign Boton[7][9] = 9'b100101000;
assign Boton[7][10] = 9'b100100100;
assign Boton[7][11] = 9'b100000100;
assign Boton[7][12] = 9'b100000100;
assign Boton[7][13] = 9'b100001001;
assign Boton[7][14] = 9'b100001001;
assign Boton[7][15] = 9'b100001001;
assign Boton[7][16] = 9'b100010010;
assign Boton[7][17] = 9'b100010111;
assign Boton[7][18] = 9'b100001101;
assign Boton[7][19] = 9'b100000100;
assign Boton[7][20] = 9'b100001001;
assign Boton[7][21] = 9'b100001001;
assign Boton[7][22] = 9'b100001001;
assign Boton[7][23] = 9'b100001001;
assign Boton[7][24] = 9'b100001001;
assign Boton[7][25] = 9'b100001001;
assign Boton[7][26] = 9'b100101001;
assign Boton[7][27] = 9'b100001001;
assign Boton[7][28] = 9'b100101001;
assign Boton[7][29] = 9'b100001001;
assign Boton[7][30] = 9'b100000101;
assign Boton[7][31] = 9'b100001001;
assign Boton[7][32] = 9'b100001001;
assign Boton[7][33] = 9'b100001001;
assign Boton[7][34] = 9'b100001001;
assign Boton[7][35] = 9'b100001001;
assign Boton[7][36] = 9'b100000100;
assign Boton[7][37] = 9'b100000100;
assign Boton[7][38] = 9'b100100100;
assign Boton[7][39] = 9'b101001000;
assign Boton[8][8] = 9'b101001000;
assign Boton[8][9] = 9'b100100100;
assign Boton[8][10] = 9'b100000100;
assign Boton[8][11] = 9'b100001001;
assign Boton[8][12] = 9'b100000100;
assign Boton[8][13] = 9'b100001001;
assign Boton[8][14] = 9'b100001001;
assign Boton[8][15] = 9'b100010011;
assign Boton[8][16] = 9'b100010111;
assign Boton[8][17] = 9'b100001101;
assign Boton[8][18] = 9'b100001001;
assign Boton[8][19] = 9'b100001001;
assign Boton[8][20] = 9'b100000101;
assign Boton[8][21] = 9'b100101001;
assign Boton[8][22] = 9'b100001001;
assign Boton[8][23] = 9'b100001001;
assign Boton[8][24] = 9'b100001001;
assign Boton[8][25] = 9'b100101001;
assign Boton[8][26] = 9'b100101001;
assign Boton[8][27] = 9'b100001001;
assign Boton[8][28] = 9'b100001001;
assign Boton[8][29] = 9'b100001001;
assign Boton[8][30] = 9'b100001001;
assign Boton[8][31] = 9'b100001001;
assign Boton[8][32] = 9'b100001001;
assign Boton[8][33] = 9'b100001001;
assign Boton[8][34] = 9'b100001001;
assign Boton[8][35] = 9'b100001001;
assign Boton[8][36] = 9'b100000100;
assign Boton[8][37] = 9'b100001001;
assign Boton[8][38] = 9'b100000100;
assign Boton[8][39] = 9'b100100000;
assign Boton[8][40] = 9'b100100100;
assign Boton[9][7] = 9'b100100100;
assign Boton[9][8] = 9'b100100100;
assign Boton[9][9] = 9'b100000000;
assign Boton[9][10] = 9'b100001101;
assign Boton[9][11] = 9'b100100100;
assign Boton[9][12] = 9'b100000100;
assign Boton[9][13] = 9'b100001001;
assign Boton[9][14] = 9'b100010111;
assign Boton[9][15] = 9'b100010011;
assign Boton[9][16] = 9'b100001101;
assign Boton[9][17] = 9'b100001001;
assign Boton[9][18] = 9'b100001001;
assign Boton[9][19] = 9'b100001001;
assign Boton[9][20] = 9'b100000101;
assign Boton[9][21] = 9'b100001001;
assign Boton[9][22] = 9'b100001001;
assign Boton[9][23] = 9'b100000101;
assign Boton[9][24] = 9'b100100101;
assign Boton[9][25] = 9'b100101001;
assign Boton[9][26] = 9'b100001001;
assign Boton[9][27] = 9'b100001001;
assign Boton[9][28] = 9'b100001001;
assign Boton[9][29] = 9'b100001001;
assign Boton[9][30] = 9'b100001001;
assign Boton[9][31] = 9'b100101001;
assign Boton[9][32] = 9'b100101001;
assign Boton[9][33] = 9'b100001001;
assign Boton[9][34] = 9'b100001001;
assign Boton[9][35] = 9'b100001001;
assign Boton[9][36] = 9'b100000100;
assign Boton[9][37] = 9'b100100100;
assign Boton[9][38] = 9'b100001101;
assign Boton[9][39] = 9'b100000100;
assign Boton[9][40] = 9'b100100100;
assign Boton[9][41] = 9'b100100100;
assign Boton[10][7] = 9'b100100100;
assign Boton[10][8] = 9'b100000000;
assign Boton[10][9] = 9'b100001101;
assign Boton[10][10] = 9'b100001001;
assign Boton[10][11] = 9'b100100000;
assign Boton[10][12] = 9'b100100100;
assign Boton[10][13] = 9'b100010010;
assign Boton[10][14] = 9'b100010111;
assign Boton[10][15] = 9'b100001101;
assign Boton[10][16] = 9'b100001001;
assign Boton[10][17] = 9'b100101001;
assign Boton[10][18] = 9'b100001001;
assign Boton[10][19] = 9'b100001001;
assign Boton[10][20] = 9'b100000100;
assign Boton[10][21] = 9'b100000100;
assign Boton[10][22] = 9'b100001001;
assign Boton[10][23] = 9'b100001101;
assign Boton[10][24] = 9'b100001101;
assign Boton[10][25] = 9'b100001101;
assign Boton[10][26] = 9'b100001101;
assign Boton[10][27] = 9'b100001001;
assign Boton[10][28] = 9'b100001001;
assign Boton[10][29] = 9'b100001001;
assign Boton[10][30] = 9'b100001001;
assign Boton[10][31] = 9'b100001001;
assign Boton[10][32] = 9'b100001001;
assign Boton[10][33] = 9'b100001001;
assign Boton[10][34] = 9'b100001001;
assign Boton[10][35] = 9'b100001001;
assign Boton[10][36] = 9'b100000100;
assign Boton[10][37] = 9'b100000000;
assign Boton[10][38] = 9'b100001001;
assign Boton[10][39] = 9'b100001101;
assign Boton[10][40] = 9'b100000000;
assign Boton[10][41] = 9'b100100100;
assign Boton[11][6] = 9'b100100100;
assign Boton[11][7] = 9'b100100000;
assign Boton[11][8] = 9'b100001001;
assign Boton[11][9] = 9'b100010010;
assign Boton[11][10] = 9'b100100100;
assign Boton[11][11] = 9'b100100000;
assign Boton[11][12] = 9'b100101000;
assign Boton[11][13] = 9'b100010011;
assign Boton[11][14] = 9'b100010010;
assign Boton[11][15] = 9'b100101001;
assign Boton[11][16] = 9'b100001001;
assign Boton[11][17] = 9'b100001001;
assign Boton[11][18] = 9'b100001001;
assign Boton[11][19] = 9'b100001001;
assign Boton[11][20] = 9'b100001001;
assign Boton[11][21] = 9'b100010010;
assign Boton[11][22] = 9'b100011111;
assign Boton[11][23] = 9'b100011111;
assign Boton[11][24] = 9'b100011111;
assign Boton[11][25] = 9'b100001101;
assign Boton[11][26] = 9'b100001001;
assign Boton[11][27] = 9'b100001001;
assign Boton[11][28] = 9'b100001101;
assign Boton[11][29] = 9'b100000100;
assign Boton[11][30] = 9'b100001001;
assign Boton[11][31] = 9'b100001001;
assign Boton[11][32] = 9'b100101001;
assign Boton[11][33] = 9'b100001001;
assign Boton[11][34] = 9'b100001001;
assign Boton[11][35] = 9'b100101001;
assign Boton[11][36] = 9'b100000100;
assign Boton[11][37] = 9'b100100000;
assign Boton[11][38] = 9'b100100100;
assign Boton[11][39] = 9'b100001101;
assign Boton[11][40] = 9'b100001001;
assign Boton[11][41] = 9'b100000000;
assign Boton[11][42] = 9'b100100100;
assign Boton[12][5] = 9'b100100100;
assign Boton[12][6] = 9'b100100100;
assign Boton[12][7] = 9'b100000100;
assign Boton[12][8] = 9'b100001101;
assign Boton[12][9] = 9'b100001001;
assign Boton[12][10] = 9'b100100100;
assign Boton[12][11] = 9'b100100000;
assign Boton[12][12] = 9'b100100100;
assign Boton[12][13] = 9'b100001101;
assign Boton[12][14] = 9'b100001101;
assign Boton[12][15] = 9'b100001001;
assign Boton[12][16] = 9'b100001001;
assign Boton[12][17] = 9'b100101001;
assign Boton[12][18] = 9'b100001001;
assign Boton[12][19] = 9'b100001001;
assign Boton[12][20] = 9'b100001001;
assign Boton[12][21] = 9'b100010111;
assign Boton[12][22] = 9'b100010111;
assign Boton[12][23] = 9'b100010111;
assign Boton[12][24] = 9'b100011111;
assign Boton[12][25] = 9'b100001110;
assign Boton[12][26] = 9'b100000100;
assign Boton[12][27] = 9'b100000000;
assign Boton[12][28] = 9'b100100100;
assign Boton[12][29] = 9'b100100100;
assign Boton[12][30] = 9'b100001001;
assign Boton[12][31] = 9'b100001001;
assign Boton[12][32] = 9'b100101001;
assign Boton[12][33] = 9'b100001001;
assign Boton[12][34] = 9'b100001001;
assign Boton[12][35] = 9'b100001001;
assign Boton[12][36] = 9'b100100100;
assign Boton[12][37] = 9'b100100100;
assign Boton[12][38] = 9'b100100000;
assign Boton[12][39] = 9'b100101001;
assign Boton[12][40] = 9'b100001110;
assign Boton[12][41] = 9'b100000100;
assign Boton[12][42] = 9'b100100000;
assign Boton[12][43] = 9'b100100100;
assign Boton[13][5] = 9'b100100100;
assign Boton[13][6] = 9'b100000000;
assign Boton[13][7] = 9'b100001001;
assign Boton[13][8] = 9'b100010010;
assign Boton[13][9] = 9'b100100100;
assign Boton[13][10] = 9'b100100100;
assign Boton[13][11] = 9'b100000000;
assign Boton[13][12] = 9'b100000000;
assign Boton[13][13] = 9'b100101000;
assign Boton[13][14] = 9'b100001001;
assign Boton[13][15] = 9'b100001001;
assign Boton[13][16] = 9'b100001001;
assign Boton[13][17] = 9'b100001001;
assign Boton[13][18] = 9'b100001001;
assign Boton[13][19] = 9'b100001001;
assign Boton[13][20] = 9'b100001101;
assign Boton[13][21] = 9'b100010111;
assign Boton[13][22] = 9'b100010111;
assign Boton[13][23] = 9'b100010111;
assign Boton[13][24] = 9'b100111111;
assign Boton[13][25] = 9'b100010010;
assign Boton[13][26] = 9'b100001001;
assign Boton[13][27] = 9'b100000000;
assign Boton[13][28] = 9'b100100000;
assign Boton[13][29] = 9'b100000100;
assign Boton[13][30] = 9'b100001001;
assign Boton[13][31] = 9'b100001001;
assign Boton[13][32] = 9'b100001001;
assign Boton[13][33] = 9'b100101001;
assign Boton[13][34] = 9'b100101001;
assign Boton[13][35] = 9'b100100100;
assign Boton[13][36] = 9'b100100100;
assign Boton[13][37] = 9'b100000000;
assign Boton[13][38] = 9'b100000000;
assign Boton[13][39] = 9'b100100100;
assign Boton[13][40] = 9'b100001101;
assign Boton[13][41] = 9'b100001101;
assign Boton[13][42] = 9'b100000000;
assign Boton[13][43] = 9'b100100100;
assign Boton[14][4] = 9'b100100100;
assign Boton[14][5] = 9'b100100000;
assign Boton[14][6] = 9'b100000100;
assign Boton[14][7] = 9'b100001101;
assign Boton[14][8] = 9'b100001101;
assign Boton[14][9] = 9'b100100000;
assign Boton[14][10] = 9'b100000000;
assign Boton[14][11] = 9'b100000000;
assign Boton[14][12] = 9'b100000000;
assign Boton[14][13] = 9'b100100100;
assign Boton[14][14] = 9'b100100100;
assign Boton[14][15] = 9'b100001001;
assign Boton[14][16] = 9'b100001001;
assign Boton[14][17] = 9'b100001001;
assign Boton[14][18] = 9'b100001001;
assign Boton[14][19] = 9'b100001101;
assign Boton[14][20] = 9'b100010011;
assign Boton[14][21] = 9'b100010111;
assign Boton[14][22] = 9'b100010111;
assign Boton[14][23] = 9'b100010111;
assign Boton[14][24] = 9'b100110111;
assign Boton[14][25] = 9'b100010010;
assign Boton[14][26] = 9'b100001001;
assign Boton[14][27] = 9'b100000000;
assign Boton[14][28] = 9'b100000000;
assign Boton[14][29] = 9'b100000100;
assign Boton[14][30] = 9'b100001001;
assign Boton[14][31] = 9'b100001001;
assign Boton[14][32] = 9'b100001001;
assign Boton[14][33] = 9'b100001001;
assign Boton[14][34] = 9'b100100100;
assign Boton[14][35] = 9'b100000000;
assign Boton[14][36] = 9'b100000000;
assign Boton[14][37] = 9'b100000000;
assign Boton[14][38] = 9'b100000000;
assign Boton[14][39] = 9'b100100000;
assign Boton[14][40] = 9'b100101101;
assign Boton[14][41] = 9'b100010010;
assign Boton[14][42] = 9'b100000100;
assign Boton[14][43] = 9'b100100000;
assign Boton[14][44] = 9'b100100100;
assign Boton[15][4] = 9'b100100100;
assign Boton[15][5] = 9'b100100000;
assign Boton[15][6] = 9'b100001001;
assign Boton[15][7] = 9'b100010010;
assign Boton[15][8] = 9'b100001001;
assign Boton[15][9] = 9'b100000000;
assign Boton[15][10] = 9'b100000000;
assign Boton[15][11] = 9'b100000000;
assign Boton[15][12] = 9'b100000000;
assign Boton[15][13] = 9'b100000000;
assign Boton[15][14] = 9'b100100100;
assign Boton[15][15] = 9'b100100100;
assign Boton[15][16] = 9'b100000101;
assign Boton[15][17] = 9'b100001001;
assign Boton[15][18] = 9'b100001001;
assign Boton[15][19] = 9'b100010011;
assign Boton[15][20] = 9'b100010111;
assign Boton[15][21] = 9'b100010111;
assign Boton[15][22] = 9'b100010111;
assign Boton[15][23] = 9'b100010111;
assign Boton[15][24] = 9'b100010111;
assign Boton[15][25] = 9'b100001101;
assign Boton[15][26] = 9'b100001001;
assign Boton[15][27] = 9'b100100100;
assign Boton[15][28] = 9'b100100000;
assign Boton[15][29] = 9'b100000100;
assign Boton[15][30] = 9'b100001101;
assign Boton[15][31] = 9'b100001001;
assign Boton[15][32] = 9'b100001001;
assign Boton[15][33] = 9'b100000100;
assign Boton[15][34] = 9'b100000000;
assign Boton[15][35] = 9'b100000000;
assign Boton[15][36] = 9'b100000000;
assign Boton[15][37] = 9'b100000000;
assign Boton[15][38] = 9'b100000000;
assign Boton[15][39] = 9'b100100000;
assign Boton[15][40] = 9'b100100100;
assign Boton[15][41] = 9'b100001110;
assign Boton[15][42] = 9'b100001001;
assign Boton[15][43] = 9'b100000000;
assign Boton[15][44] = 9'b100100100;
assign Boton[16][4] = 9'b100100000;
assign Boton[16][5] = 9'b100000100;
assign Boton[16][6] = 9'b100001101;
assign Boton[16][7] = 9'b100001110;
assign Boton[16][8] = 9'b100100100;
assign Boton[16][9] = 9'b100000000;
assign Boton[16][10] = 9'b100000000;
assign Boton[16][11] = 9'b100000000;
assign Boton[16][12] = 9'b100000000;
assign Boton[16][13] = 9'b100100100;
assign Boton[16][14] = 9'b100100100;
assign Boton[16][15] = 9'b100100000;
assign Boton[16][16] = 9'b100100100;
assign Boton[16][17] = 9'b100100000;
assign Boton[16][18] = 9'b100101001;
assign Boton[16][19] = 9'b100010111;
assign Boton[16][20] = 9'b100010011;
assign Boton[16][21] = 9'b100010011;
assign Boton[16][22] = 9'b100010011;
assign Boton[16][23] = 9'b100010011;
assign Boton[16][24] = 9'b100001101;
assign Boton[16][25] = 9'b100001001;
assign Boton[16][26] = 9'b100000101;
assign Boton[16][27] = 9'b100000000;
assign Boton[16][28] = 9'b100000000;
assign Boton[16][29] = 9'b100000100;
assign Boton[16][30] = 9'b100001101;
assign Boton[16][31] = 9'b100100100;
assign Boton[16][32] = 9'b100100100;
assign Boton[16][33] = 9'b100100100;
assign Boton[16][34] = 9'b100100000;
assign Boton[16][35] = 9'b100100100;
assign Boton[16][36] = 9'b100100100;
assign Boton[16][37] = 9'b100100100;
assign Boton[16][38] = 9'b100100100;
assign Boton[16][39] = 9'b100000000;
assign Boton[16][40] = 9'b100000000;
assign Boton[16][41] = 9'b100001101;
assign Boton[16][42] = 9'b100001101;
assign Boton[16][43] = 9'b100000100;
assign Boton[16][44] = 9'b100100000;
assign Boton[16][45] = 9'b100100100;
assign Boton[17][3] = 9'b100100100;
assign Boton[17][4] = 9'b100100000;
assign Boton[17][5] = 9'b100000100;
assign Boton[17][6] = 9'b100001101;
assign Boton[17][7] = 9'b100001101;
assign Boton[17][8] = 9'b100000000;
assign Boton[17][9] = 9'b100100100;
assign Boton[17][10] = 9'b100100100;
assign Boton[17][11] = 9'b100100100;
assign Boton[17][12] = 9'b100100000;
assign Boton[17][13] = 9'b100000000;
assign Boton[17][14] = 9'b100000100;
assign Boton[17][15] = 9'b100100100;
assign Boton[17][16] = 9'b100100100;
assign Boton[17][17] = 9'b100000000;
assign Boton[17][18] = 9'b100001001;
assign Boton[17][19] = 9'b100011111;
assign Boton[17][20] = 9'b100001101;
assign Boton[17][21] = 9'b100001001;
assign Boton[17][22] = 9'b100001001;
assign Boton[17][23] = 9'b100001001;
assign Boton[17][24] = 9'b100001001;
assign Boton[17][25] = 9'b100000101;
assign Boton[17][26] = 9'b100100100;
assign Boton[17][27] = 9'b100000000;
assign Boton[17][28] = 9'b100000000;
assign Boton[17][29] = 9'b100000100;
assign Boton[17][30] = 9'b100001101;
assign Boton[17][31] = 9'b100000000;
assign Boton[17][32] = 9'b100000000;
assign Boton[17][33] = 9'b100000100;
assign Boton[17][34] = 9'b100000100;
assign Boton[17][35] = 9'b100000000;
assign Boton[17][36] = 9'b100000000;
assign Boton[17][37] = 9'b100000000;
assign Boton[17][38] = 9'b100100100;
assign Boton[17][39] = 9'b100100100;
assign Boton[17][40] = 9'b100100000;
assign Boton[17][41] = 9'b100001001;
assign Boton[17][42] = 9'b100001110;
assign Boton[17][43] = 9'b100001001;
assign Boton[17][44] = 9'b100100000;
assign Boton[17][45] = 9'b100100100;
assign Boton[18][3] = 9'b100100100;
assign Boton[18][4] = 9'b100100000;
assign Boton[18][5] = 9'b100001001;
assign Boton[18][6] = 9'b100001110;
assign Boton[18][7] = 9'b100001001;
assign Boton[18][8] = 9'b100000000;
assign Boton[18][9] = 9'b100100100;
assign Boton[18][10] = 9'b100100100;
assign Boton[18][11] = 9'b100100100;
assign Boton[18][12] = 9'b100000100;
assign Boton[18][13] = 9'b100001001;
assign Boton[18][14] = 9'b100000101;
assign Boton[18][15] = 9'b100100100;
assign Boton[18][16] = 9'b100000000;
assign Boton[18][17] = 9'b100100000;
assign Boton[18][18] = 9'b100001001;
assign Boton[18][19] = 9'b100010111;
assign Boton[18][20] = 9'b100001001;
assign Boton[18][21] = 9'b100000100;
assign Boton[18][22] = 9'b100100100;
assign Boton[18][23] = 9'b100100100;
assign Boton[18][24] = 9'b100000100;
assign Boton[18][25] = 9'b100000000;
assign Boton[18][26] = 9'b100000000;
assign Boton[18][27] = 9'b100100100;
assign Boton[18][28] = 9'b100000000;
assign Boton[18][29] = 9'b100001001;
assign Boton[18][30] = 9'b100001101;
assign Boton[18][31] = 9'b100000000;
assign Boton[18][32] = 9'b100100100;
assign Boton[18][33] = 9'b100100000;
assign Boton[18][34] = 9'b100000101;
assign Boton[18][35] = 9'b100000101;
assign Boton[18][36] = 9'b100000000;
assign Boton[18][37] = 9'b100100000;
assign Boton[18][38] = 9'b100100100;
assign Boton[18][39] = 9'b100000000;
assign Boton[18][40] = 9'b100100000;
assign Boton[18][41] = 9'b100101001;
assign Boton[18][42] = 9'b100001110;
assign Boton[18][43] = 9'b100001001;
assign Boton[18][44] = 9'b100000000;
assign Boton[18][45] = 9'b100100100;
assign Boton[19][3] = 9'b100100000;
assign Boton[19][4] = 9'b100100100;
assign Boton[19][5] = 9'b100001101;
assign Boton[19][6] = 9'b100010010;
assign Boton[19][7] = 9'b100000100;
assign Boton[19][8] = 9'b100100000;
assign Boton[19][9] = 9'b100100000;
assign Boton[19][10] = 9'b100000000;
assign Boton[19][11] = 9'b100000100;
assign Boton[19][12] = 9'b100001001;
assign Boton[19][13] = 9'b100001001;
assign Boton[19][14] = 9'b100000100;
assign Boton[19][15] = 9'b100100100;
assign Boton[19][16] = 9'b100100100;
assign Boton[19][17] = 9'b100100100;
assign Boton[19][18] = 9'b100001101;
assign Boton[19][19] = 9'b100010111;
assign Boton[19][20] = 9'b100010010;
assign Boton[19][21] = 9'b100001001;
assign Boton[19][22] = 9'b100000000;
assign Boton[19][23] = 9'b100100000;
assign Boton[19][24] = 9'b100000000;
assign Boton[19][25] = 9'b100000000;
assign Boton[19][26] = 9'b100100100;
assign Boton[19][27] = 9'b100000000;
assign Boton[19][28] = 9'b100001101;
assign Boton[19][29] = 9'b100001110;
assign Boton[19][30] = 9'b100001101;
assign Boton[19][31] = 9'b100100100;
assign Boton[19][32] = 9'b100000000;
assign Boton[19][33] = 9'b100000000;
assign Boton[19][34] = 9'b100000100;
assign Boton[19][35] = 9'b100001001;
assign Boton[19][36] = 9'b100001001;
assign Boton[19][37] = 9'b100000100;
assign Boton[19][38] = 9'b100000000;
assign Boton[19][39] = 9'b100100100;
assign Boton[19][40] = 9'b100000000;
assign Boton[19][41] = 9'b100100100;
assign Boton[19][42] = 9'b100010010;
assign Boton[19][43] = 9'b100001101;
assign Boton[19][44] = 9'b100000100;
assign Boton[19][45] = 9'b100100100;
assign Boton[20][3] = 9'b100000000;
assign Boton[20][4] = 9'b100000100;
assign Boton[20][5] = 9'b100001101;
assign Boton[20][6] = 9'b100001101;
assign Boton[20][7] = 9'b100000100;
assign Boton[20][8] = 9'b100100000;
assign Boton[20][9] = 9'b100000000;
assign Boton[20][10] = 9'b100000100;
assign Boton[20][11] = 9'b100001001;
assign Boton[20][12] = 9'b100001001;
assign Boton[20][13] = 9'b100101001;
assign Boton[20][14] = 9'b100000100;
assign Boton[20][15] = 9'b100100000;
assign Boton[20][16] = 9'b100100100;
assign Boton[20][17] = 9'b100100000;
assign Boton[20][18] = 9'b100001101;
assign Boton[20][19] = 9'b100010011;
assign Boton[20][20] = 9'b100101000;
assign Boton[20][21] = 9'b100001101;
assign Boton[20][22] = 9'b100001101;
assign Boton[20][23] = 9'b100000000;
assign Boton[20][24] = 9'b100000000;
assign Boton[20][25] = 9'b100000000;
assign Boton[20][26] = 9'b100000100;
assign Boton[20][27] = 9'b100001001;
assign Boton[20][28] = 9'b100001101;
assign Boton[20][29] = 9'b100001101;
assign Boton[20][30] = 9'b100001101;
assign Boton[20][31] = 9'b100100100;
assign Boton[20][32] = 9'b100100000;
assign Boton[20][33] = 9'b100100000;
assign Boton[20][34] = 9'b100000100;
assign Boton[20][35] = 9'b100001001;
assign Boton[20][36] = 9'b100001001;
assign Boton[20][37] = 9'b100001001;
assign Boton[20][38] = 9'b100000100;
assign Boton[20][39] = 9'b100000000;
assign Boton[20][40] = 9'b100100000;
assign Boton[20][41] = 9'b100100100;
assign Boton[20][42] = 9'b100010010;
assign Boton[20][43] = 9'b100001101;
assign Boton[20][44] = 9'b100000100;
assign Boton[20][45] = 9'b100100000;
assign Boton[20][46] = 9'b100100100;
assign Boton[21][2] = 9'b100100100;
assign Boton[21][3] = 9'b100100000;
assign Boton[21][4] = 9'b100001001;
assign Boton[21][5] = 9'b100001101;
assign Boton[21][6] = 9'b100001101;
assign Boton[21][7] = 9'b100100000;
assign Boton[21][8] = 9'b100000000;
assign Boton[21][9] = 9'b100000100;
assign Boton[21][10] = 9'b100101001;
assign Boton[21][11] = 9'b100001001;
assign Boton[21][12] = 9'b100001001;
assign Boton[21][13] = 9'b100001001;
assign Boton[21][14] = 9'b100001001;
assign Boton[21][15] = 9'b100000000;
assign Boton[21][16] = 9'b100100000;
assign Boton[21][17] = 9'b100100000;
assign Boton[21][18] = 9'b100001101;
assign Boton[21][19] = 9'b100001101;
assign Boton[21][20] = 9'b100100000;
assign Boton[21][21] = 9'b100100100;
assign Boton[21][22] = 9'b100001101;
assign Boton[21][23] = 9'b100001001;
assign Boton[21][24] = 9'b100000100;
assign Boton[21][25] = 9'b100000000;
assign Boton[21][26] = 9'b100001101;
assign Boton[21][27] = 9'b100101101;
assign Boton[21][28] = 9'b100100100;
assign Boton[21][29] = 9'b100000100;
assign Boton[21][30] = 9'b100001101;
assign Boton[21][31] = 9'b100100100;
assign Boton[21][32] = 9'b100100000;
assign Boton[21][33] = 9'b100000100;
assign Boton[21][34] = 9'b100101001;
assign Boton[21][35] = 9'b100101001;
assign Boton[21][36] = 9'b100101001;
assign Boton[21][37] = 9'b100001001;
assign Boton[21][38] = 9'b100001001;
assign Boton[21][39] = 9'b100000100;
assign Boton[21][40] = 9'b100000000;
assign Boton[21][41] = 9'b100100100;
assign Boton[21][42] = 9'b100001101;
assign Boton[21][43] = 9'b100001110;
assign Boton[21][44] = 9'b100001001;
assign Boton[21][45] = 9'b100100100;
assign Boton[21][46] = 9'b100100100;
assign Boton[22][2] = 9'b100100100;
assign Boton[22][3] = 9'b100100100;
assign Boton[22][4] = 9'b100001001;
assign Boton[22][5] = 9'b100001101;
assign Boton[22][6] = 9'b100001101;
assign Boton[22][7] = 9'b100000000;
assign Boton[22][8] = 9'b100000100;
assign Boton[22][9] = 9'b100101001;
assign Boton[22][10] = 9'b100101001;
assign Boton[22][11] = 9'b100101001;
assign Boton[22][12] = 9'b100101001;
assign Boton[22][13] = 9'b100001001;
assign Boton[22][14] = 9'b100001001;
assign Boton[22][15] = 9'b100001001;
assign Boton[22][16] = 9'b100000000;
assign Boton[22][17] = 9'b100100000;
assign Boton[22][18] = 9'b100001101;
assign Boton[22][19] = 9'b100010011;
assign Boton[22][20] = 9'b100101001;
assign Boton[22][21] = 9'b110010001;
assign Boton[22][22] = 9'b101001001;
assign Boton[22][23] = 9'b100001001;
assign Boton[22][24] = 9'b100000100;
assign Boton[22][25] = 9'b100000100;
assign Boton[22][26] = 9'b100101001;
assign Boton[22][27] = 9'b110010001;
assign Boton[22][28] = 9'b101001000;
assign Boton[22][29] = 9'b100000100;
assign Boton[22][30] = 9'b100001101;
assign Boton[22][31] = 9'b100000000;
assign Boton[22][32] = 9'b100000000;
assign Boton[22][33] = 9'b100001001;
assign Boton[22][34] = 9'b100101001;
assign Boton[22][35] = 9'b100001001;
assign Boton[22][36] = 9'b100101001;
assign Boton[22][37] = 9'b100001001;
assign Boton[22][38] = 9'b100001001;
assign Boton[22][39] = 9'b100001001;
assign Boton[22][40] = 9'b100000100;
assign Boton[22][41] = 9'b100100000;
assign Boton[22][42] = 9'b100001101;
assign Boton[22][43] = 9'b100001110;
assign Boton[22][44] = 9'b100001001;
assign Boton[22][45] = 9'b100100000;
assign Boton[22][46] = 9'b100100100;
assign Boton[23][2] = 9'b100100100;
assign Boton[23][3] = 9'b100100000;
assign Boton[23][4] = 9'b100001001;
assign Boton[23][5] = 9'b100001101;
assign Boton[23][6] = 9'b100001101;
assign Boton[23][7] = 9'b100000000;
assign Boton[23][8] = 9'b100001001;
assign Boton[23][9] = 9'b100001001;
assign Boton[23][10] = 9'b100001001;
assign Boton[23][11] = 9'b100001001;
assign Boton[23][12] = 9'b100001001;
assign Boton[23][13] = 9'b100001001;
assign Boton[23][14] = 9'b100101001;
assign Boton[23][15] = 9'b100101001;
assign Boton[23][16] = 9'b100001001;
assign Boton[23][17] = 9'b100000000;
assign Boton[23][18] = 9'b100001001;
assign Boton[23][19] = 9'b100010111;
assign Boton[23][20] = 9'b100001101;
assign Boton[23][21] = 9'b100001001;
assign Boton[23][22] = 9'b100100100;
assign Boton[23][23] = 9'b100000100;
assign Boton[23][24] = 9'b100000100;
assign Boton[23][25] = 9'b100000100;
assign Boton[23][26] = 9'b100100100;
assign Boton[23][27] = 9'b100100100;
assign Boton[23][28] = 9'b100000100;
assign Boton[23][29] = 9'b100001001;
assign Boton[23][30] = 9'b100001101;
assign Boton[23][31] = 9'b100000000;
assign Boton[23][32] = 9'b100001001;
assign Boton[23][33] = 9'b100001001;
assign Boton[23][34] = 9'b100101001;
assign Boton[23][35] = 9'b100101001;
assign Boton[23][36] = 9'b100101001;
assign Boton[23][37] = 9'b100101001;
assign Boton[23][38] = 9'b100101001;
assign Boton[23][39] = 9'b100101001;
assign Boton[23][40] = 9'b100001001;
assign Boton[23][41] = 9'b100000000;
assign Boton[23][42] = 9'b100001001;
assign Boton[23][43] = 9'b100001110;
assign Boton[23][44] = 9'b100001001;
assign Boton[23][45] = 9'b100100100;
assign Boton[23][46] = 9'b100100100;
assign Boton[24][2] = 9'b100100100;
assign Boton[24][3] = 9'b100100000;
assign Boton[24][4] = 9'b100001001;
assign Boton[24][5] = 9'b100001110;
assign Boton[24][6] = 9'b100001101;
assign Boton[24][7] = 9'b100000100;
assign Boton[24][8] = 9'b100001001;
assign Boton[24][9] = 9'b100001001;
assign Boton[24][10] = 9'b100001001;
assign Boton[24][11] = 9'b100001001;
assign Boton[24][12] = 9'b100001001;
assign Boton[24][13] = 9'b100001001;
assign Boton[24][14] = 9'b100001001;
assign Boton[24][15] = 9'b100101001;
assign Boton[24][16] = 9'b100001001;
assign Boton[24][17] = 9'b100001001;
assign Boton[24][18] = 9'b100000100;
assign Boton[24][19] = 9'b100010011;
assign Boton[24][20] = 9'b100001101;
assign Boton[24][21] = 9'b100001001;
assign Boton[24][22] = 9'b100000100;
assign Boton[24][23] = 9'b100000100;
assign Boton[24][24] = 9'b100001001;
assign Boton[24][25] = 9'b100000101;
assign Boton[24][26] = 9'b100000000;
assign Boton[24][27] = 9'b100000000;
assign Boton[24][28] = 9'b100000000;
assign Boton[24][29] = 9'b100001001;
assign Boton[24][30] = 9'b100001101;
assign Boton[24][31] = 9'b100001001;
assign Boton[24][32] = 9'b100101001;
assign Boton[24][33] = 9'b100001001;
assign Boton[24][34] = 9'b100001001;
assign Boton[24][35] = 9'b100101001;
assign Boton[24][36] = 9'b100001001;
assign Boton[24][37] = 9'b100101001;
assign Boton[24][38] = 9'b100101001;
assign Boton[24][39] = 9'b100001001;
assign Boton[24][40] = 9'b100001001;
assign Boton[24][41] = 9'b100000100;
assign Boton[24][42] = 9'b100001001;
assign Boton[24][43] = 9'b100001110;
assign Boton[24][44] = 9'b100001001;
assign Boton[24][45] = 9'b100100000;
assign Boton[24][46] = 9'b100100100;
assign Boton[25][2] = 9'b100100100;
assign Boton[25][3] = 9'b100100000;
assign Boton[25][4] = 9'b100001001;
assign Boton[25][5] = 9'b100001110;
assign Boton[25][6] = 9'b100001101;
assign Boton[25][7] = 9'b100000101;
assign Boton[25][8] = 9'b100101001;
assign Boton[25][9] = 9'b100101001;
assign Boton[25][10] = 9'b100101001;
assign Boton[25][11] = 9'b100001001;
assign Boton[25][12] = 9'b100001001;
assign Boton[25][13] = 9'b100001001;
assign Boton[25][14] = 9'b100101001;
assign Boton[25][15] = 9'b100101001;
assign Boton[25][16] = 9'b100101001;
assign Boton[25][17] = 9'b100001001;
assign Boton[25][18] = 9'b100001001;
assign Boton[25][19] = 9'b100110010;
assign Boton[25][20] = 9'b110010001;
assign Boton[25][21] = 9'b100101001;
assign Boton[25][22] = 9'b100000000;
assign Boton[25][23] = 9'b100000101;
assign Boton[25][24] = 9'b100001001;
assign Boton[25][25] = 9'b100001001;
assign Boton[25][26] = 9'b100000100;
assign Boton[25][27] = 9'b100000000;
assign Boton[25][28] = 9'b101001000;
assign Boton[25][29] = 9'b101001101;
assign Boton[25][30] = 9'b100001101;
assign Boton[25][31] = 9'b100001001;
assign Boton[25][32] = 9'b100001001;
assign Boton[25][33] = 9'b100101001;
assign Boton[25][34] = 9'b100101001;
assign Boton[25][35] = 9'b100101001;
assign Boton[25][36] = 9'b100101001;
assign Boton[25][37] = 9'b100001001;
assign Boton[25][38] = 9'b100001001;
assign Boton[25][39] = 9'b100001001;
assign Boton[25][40] = 9'b100001001;
assign Boton[25][41] = 9'b100000101;
assign Boton[25][42] = 9'b100001001;
assign Boton[25][43] = 9'b100001110;
assign Boton[25][44] = 9'b100001001;
assign Boton[25][45] = 9'b100000000;
assign Boton[25][46] = 9'b100100100;
assign Boton[26][2] = 9'b100000000;
assign Boton[26][3] = 9'b100100000;
assign Boton[26][4] = 9'b100001001;
assign Boton[26][5] = 9'b100001101;
assign Boton[26][6] = 9'b100010010;
assign Boton[26][7] = 9'b100001001;
assign Boton[26][8] = 9'b100001001;
assign Boton[26][9] = 9'b100101001;
assign Boton[26][10] = 9'b100101001;
assign Boton[26][11] = 9'b100101001;
assign Boton[26][12] = 9'b100101001;
assign Boton[26][13] = 9'b100101001;
assign Boton[26][14] = 9'b100101001;
assign Boton[26][15] = 9'b100101001;
assign Boton[26][16] = 9'b100101001;
assign Boton[26][17] = 9'b100101001;
assign Boton[26][18] = 9'b100001001;
assign Boton[26][19] = 9'b100010010;
assign Boton[26][20] = 9'b111110110;
assign Boton[26][21] = 9'b111110110;
assign Boton[26][22] = 9'b101101001;
assign Boton[26][23] = 9'b100001001;
assign Boton[26][24] = 9'b100000100;
assign Boton[26][25] = 9'b100000100;
assign Boton[26][26] = 9'b100101001;
assign Boton[26][27] = 9'b110001101;
assign Boton[26][28] = 9'b111110101;
assign Boton[26][29] = 9'b101101101;
assign Boton[26][30] = 9'b100001101;
assign Boton[26][31] = 9'b100001001;
assign Boton[26][32] = 9'b100001001;
assign Boton[26][33] = 9'b100001001;
assign Boton[26][34] = 9'b100001001;
assign Boton[26][35] = 9'b100001001;
assign Boton[26][36] = 9'b100001001;
assign Boton[26][37] = 9'b100001001;
assign Boton[26][38] = 9'b100001001;
assign Boton[26][39] = 9'b100001001;
assign Boton[26][40] = 9'b100001001;
assign Boton[26][41] = 9'b100001001;
assign Boton[26][42] = 9'b100001101;
assign Boton[26][43] = 9'b100001110;
assign Boton[26][44] = 9'b100001001;
assign Boton[26][45] = 9'b100000000;
assign Boton[26][46] = 9'b100100100;
assign Boton[27][2] = 9'b100000000;
assign Boton[27][3] = 9'b100000000;
assign Boton[27][4] = 9'b100001001;
assign Boton[27][5] = 9'b100001110;
assign Boton[27][6] = 9'b100010010;
assign Boton[27][7] = 9'b100001001;
assign Boton[27][8] = 9'b100101001;
assign Boton[27][9] = 9'b100101001;
assign Boton[27][10] = 9'b100101001;
assign Boton[27][11] = 9'b100001001;
assign Boton[27][12] = 9'b100001001;
assign Boton[27][13] = 9'b100001001;
assign Boton[27][14] = 9'b100001001;
assign Boton[27][15] = 9'b100101001;
assign Boton[27][16] = 9'b100101001;
assign Boton[27][17] = 9'b100001001;
assign Boton[27][18] = 9'b100001001;
assign Boton[27][19] = 9'b100010010;
assign Boton[27][20] = 9'b110110010;
assign Boton[27][21] = 9'b111110110;
assign Boton[27][22] = 9'b111111110;
assign Boton[27][23] = 9'b110110010;
assign Boton[27][24] = 9'b100101001;
assign Boton[27][25] = 9'b100101001;
assign Boton[27][26] = 9'b111110110;
assign Boton[27][27] = 9'b111110110;
assign Boton[27][28] = 9'b110110001;
assign Boton[27][29] = 9'b101001101;
assign Boton[27][30] = 9'b100001001;
assign Boton[27][31] = 9'b100001001;
assign Boton[27][32] = 9'b100001001;
assign Boton[27][33] = 9'b100001001;
assign Boton[27][34] = 9'b100001001;
assign Boton[27][35] = 9'b100101001;
assign Boton[27][36] = 9'b100001001;
assign Boton[27][37] = 9'b100001001;
assign Boton[27][38] = 9'b100101001;
assign Boton[27][39] = 9'b100101001;
assign Boton[27][40] = 9'b100101001;
assign Boton[27][41] = 9'b100101001;
assign Boton[27][42] = 9'b100001110;
assign Boton[27][43] = 9'b100001110;
assign Boton[27][44] = 9'b100001001;
assign Boton[27][45] = 9'b100100000;
assign Boton[27][46] = 9'b100100100;
assign Boton[28][2] = 9'b100000100;
assign Boton[28][3] = 9'b100100000;
assign Boton[28][4] = 9'b100001001;
assign Boton[28][5] = 9'b100001110;
assign Boton[28][6] = 9'b100010010;
assign Boton[28][7] = 9'b100001001;
assign Boton[28][8] = 9'b100101001;
assign Boton[28][9] = 9'b100001001;
assign Boton[28][10] = 9'b100001001;
assign Boton[28][11] = 9'b100001001;
assign Boton[28][12] = 9'b100001001;
assign Boton[28][13] = 9'b100001001;
assign Boton[28][14] = 9'b100001001;
assign Boton[28][15] = 9'b100101001;
assign Boton[28][16] = 9'b100001001;
assign Boton[28][17] = 9'b100001001;
assign Boton[28][18] = 9'b100001001;
assign Boton[28][19] = 9'b100001101;
assign Boton[28][20] = 9'b110010010;
assign Boton[28][21] = 9'b111111110;
assign Boton[28][22] = 9'b110110010;
assign Boton[28][23] = 9'b110010001;
assign Boton[28][24] = 9'b110010001;
assign Boton[28][25] = 9'b110010001;
assign Boton[28][26] = 9'b110010001;
assign Boton[28][27] = 9'b110110010;
assign Boton[28][28] = 9'b111110001;
assign Boton[28][29] = 9'b101001101;
assign Boton[28][30] = 9'b100001001;
assign Boton[28][31] = 9'b100101001;
assign Boton[28][32] = 9'b100101001;
assign Boton[28][33] = 9'b100101001;
assign Boton[28][34] = 9'b100001001;
assign Boton[28][35] = 9'b100001001;
assign Boton[28][36] = 9'b100001001;
assign Boton[28][37] = 9'b100101001;
assign Boton[28][38] = 9'b100101001;
assign Boton[28][39] = 9'b100101001;
assign Boton[28][40] = 9'b100101001;
assign Boton[28][41] = 9'b100001001;
assign Boton[28][42] = 9'b100010010;
assign Boton[28][43] = 9'b100010010;
assign Boton[28][44] = 9'b100001001;
assign Boton[28][45] = 9'b100100000;
assign Boton[28][46] = 9'b100100100;
assign Boton[29][3] = 9'b100100100;
assign Boton[29][4] = 9'b100100100;
assign Boton[29][5] = 9'b100001101;
assign Boton[29][6] = 9'b100010010;
assign Boton[29][7] = 9'b100001001;
assign Boton[29][8] = 9'b100101001;
assign Boton[29][9] = 9'b100001001;
assign Boton[29][10] = 9'b100101001;
assign Boton[29][11] = 9'b100101001;
assign Boton[29][12] = 9'b100101001;
assign Boton[29][13] = 9'b100101001;
assign Boton[29][14] = 9'b100001001;
assign Boton[29][15] = 9'b100001001;
assign Boton[29][16] = 9'b100001001;
assign Boton[29][17] = 9'b100001001;
assign Boton[29][18] = 9'b100001001;
assign Boton[29][19] = 9'b100001001;
assign Boton[29][20] = 9'b110010110;
assign Boton[29][21] = 9'b111110010;
assign Boton[29][22] = 9'b101001000;
assign Boton[29][23] = 9'b101001001;
assign Boton[29][24] = 9'b101101101;
assign Boton[29][25] = 9'b101101101;
assign Boton[29][26] = 9'b100100100;
assign Boton[29][27] = 9'b101101101;
assign Boton[29][28] = 9'b111110001;
assign Boton[29][29] = 9'b100101101;
assign Boton[29][30] = 9'b100001001;
assign Boton[29][31] = 9'b100001001;
assign Boton[29][32] = 9'b100101001;
assign Boton[29][33] = 9'b100101001;
assign Boton[29][34] = 9'b100101001;
assign Boton[29][35] = 9'b100001001;
assign Boton[29][36] = 9'b100001001;
assign Boton[29][37] = 9'b100101001;
assign Boton[29][38] = 9'b100001001;
assign Boton[29][39] = 9'b100001001;
assign Boton[29][40] = 9'b100001001;
assign Boton[29][41] = 9'b100001001;
assign Boton[29][42] = 9'b100010010;
assign Boton[29][43] = 9'b100001110;
assign Boton[29][44] = 9'b100000100;
assign Boton[29][45] = 9'b100100000;
assign Boton[30][3] = 9'b100000000;
assign Boton[30][4] = 9'b100100100;
assign Boton[30][5] = 9'b100001101;
assign Boton[30][6] = 9'b100010011;
assign Boton[30][7] = 9'b100001101;
assign Boton[30][8] = 9'b100101001;
assign Boton[30][9] = 9'b100001001;
assign Boton[30][10] = 9'b100001001;
assign Boton[30][11] = 9'b100101001;
assign Boton[30][12] = 9'b100101001;
assign Boton[30][13] = 9'b100001001;
assign Boton[30][14] = 9'b100001001;
assign Boton[30][15] = 9'b100101001;
assign Boton[30][16] = 9'b100001001;
assign Boton[30][17] = 9'b100001001;
assign Boton[30][18] = 9'b100001001;
assign Boton[30][19] = 9'b100000100;
assign Boton[30][20] = 9'b101110001;
assign Boton[30][21] = 9'b111110110;
assign Boton[30][22] = 9'b110010001;
assign Boton[30][23] = 9'b101101101;
assign Boton[30][24] = 9'b101101101;
assign Boton[30][25] = 9'b101101101;
assign Boton[30][26] = 9'b101101101;
assign Boton[30][27] = 9'b110110001;
assign Boton[30][28] = 9'b110110010;
assign Boton[30][29] = 9'b100001101;
assign Boton[30][30] = 9'b100001001;
assign Boton[30][31] = 9'b100001001;
assign Boton[30][32] = 9'b100001001;
assign Boton[30][33] = 9'b100001001;
assign Boton[30][34] = 9'b100101001;
assign Boton[30][35] = 9'b100001001;
assign Boton[30][36] = 9'b100001001;
assign Boton[30][37] = 9'b100001001;
assign Boton[30][38] = 9'b100001001;
assign Boton[30][39] = 9'b100101001;
assign Boton[30][40] = 9'b100001001;
assign Boton[30][41] = 9'b100001001;
assign Boton[30][42] = 9'b100010010;
assign Boton[30][43] = 9'b100001101;
assign Boton[30][44] = 9'b100000100;
assign Boton[30][45] = 9'b100100100;
assign Boton[31][3] = 9'b100000000;
assign Boton[31][4] = 9'b100100000;
assign Boton[31][5] = 9'b100001001;
assign Boton[31][6] = 9'b100010011;
assign Boton[31][7] = 9'b100001110;
assign Boton[31][8] = 9'b100001001;
assign Boton[31][9] = 9'b100001001;
assign Boton[31][10] = 9'b100001001;
assign Boton[31][11] = 9'b100001001;
assign Boton[31][12] = 9'b100001001;
assign Boton[31][13] = 9'b100001001;
assign Boton[31][14] = 9'b100101001;
assign Boton[31][15] = 9'b100101001;
assign Boton[31][16] = 9'b100101001;
assign Boton[31][17] = 9'b100001001;
assign Boton[31][18] = 9'b100001001;
assign Boton[31][19] = 9'b100001001;
assign Boton[31][20] = 9'b100100100;
assign Boton[31][21] = 9'b111110110;
assign Boton[31][22] = 9'b111110110;
assign Boton[31][23] = 9'b111110110;
assign Boton[31][24] = 9'b111111110;
assign Boton[31][25] = 9'b111110010;
assign Boton[31][26] = 9'b110010001;
assign Boton[31][27] = 9'b111110110;
assign Boton[31][28] = 9'b110010001;
assign Boton[31][29] = 9'b100000100;
assign Boton[31][30] = 9'b100001001;
assign Boton[31][31] = 9'b100001001;
assign Boton[31][32] = 9'b100101001;
assign Boton[31][33] = 9'b100101001;
assign Boton[31][34] = 9'b100101001;
assign Boton[31][35] = 9'b100101001;
assign Boton[31][36] = 9'b100001001;
assign Boton[31][37] = 9'b100001001;
assign Boton[31][38] = 9'b100001001;
assign Boton[31][39] = 9'b100101001;
assign Boton[31][40] = 9'b100101001;
assign Boton[31][41] = 9'b100001101;
assign Boton[31][42] = 9'b100010011;
assign Boton[31][43] = 9'b100001101;
assign Boton[31][44] = 9'b100100100;
assign Boton[31][45] = 9'b100100100;
assign Boton[32][3] = 9'b100000000;
assign Boton[32][4] = 9'b100000000;
assign Boton[32][5] = 9'b100100100;
assign Boton[32][6] = 9'b100010010;
assign Boton[32][7] = 9'b100010011;
assign Boton[32][8] = 9'b100001001;
assign Boton[32][9] = 9'b100101001;
assign Boton[32][10] = 9'b100001001;
assign Boton[32][11] = 9'b100001001;
assign Boton[32][12] = 9'b100100100;
assign Boton[32][13] = 9'b100100100;
assign Boton[32][14] = 9'b100100100;
assign Boton[32][15] = 9'b100100101;
assign Boton[32][16] = 9'b100001001;
assign Boton[32][17] = 9'b100001001;
assign Boton[32][18] = 9'b100001001;
assign Boton[32][19] = 9'b100001001;
assign Boton[32][20] = 9'b100000101;
assign Boton[32][21] = 9'b110001101;
assign Boton[32][22] = 9'b111110110;
assign Boton[32][23] = 9'b101101101;
assign Boton[32][24] = 9'b101101101;
assign Boton[32][25] = 9'b101101101;
assign Boton[32][26] = 9'b101101101;
assign Boton[32][27] = 9'b111110110;
assign Boton[32][28] = 9'b101001000;
assign Boton[32][29] = 9'b100000100;
assign Boton[32][30] = 9'b100101001;
assign Boton[32][31] = 9'b100001001;
assign Boton[32][32] = 9'b100101001;
assign Boton[32][33] = 9'b100100100;
assign Boton[32][34] = 9'b100100100;
assign Boton[32][35] = 9'b100100100;
assign Boton[32][36] = 9'b100101001;
assign Boton[32][37] = 9'b100001001;
assign Boton[32][38] = 9'b100101001;
assign Boton[32][39] = 9'b100001001;
assign Boton[32][40] = 9'b100001001;
assign Boton[32][41] = 9'b100010010;
assign Boton[32][42] = 9'b100010111;
assign Boton[32][43] = 9'b100001001;
assign Boton[32][44] = 9'b100100000;
assign Boton[32][45] = 9'b100100100;
assign Boton[33][4] = 9'b100000000;
assign Boton[33][5] = 9'b100100100;
assign Boton[33][6] = 9'b100001101;
assign Boton[33][7] = 9'b100010111;
assign Boton[33][8] = 9'b100001001;
assign Boton[33][9] = 9'b100001001;
assign Boton[33][10] = 9'b100001001;
assign Boton[33][11] = 9'b100100100;
assign Boton[33][12] = 9'b100100000;
assign Boton[33][13] = 9'b100100100;
assign Boton[33][14] = 9'b100100100;
assign Boton[33][15] = 9'b100100000;
assign Boton[33][16] = 9'b100100100;
assign Boton[33][17] = 9'b100100100;
assign Boton[33][18] = 9'b100101001;
assign Boton[33][19] = 9'b100001001;
assign Boton[33][20] = 9'b100001001;
assign Boton[33][21] = 9'b100000100;
assign Boton[33][22] = 9'b110010001;
assign Boton[33][23] = 9'b111111110;
assign Boton[33][24] = 9'b111110110;
assign Boton[33][25] = 9'b111111110;
assign Boton[33][26] = 9'b111110110;
assign Boton[33][27] = 9'b101101001;
assign Boton[33][28] = 9'b100000100;
assign Boton[33][29] = 9'b100001001;
assign Boton[33][30] = 9'b100000101;
assign Boton[33][31] = 9'b100100100;
assign Boton[33][32] = 9'b100100100;
assign Boton[33][33] = 9'b100000000;
assign Boton[33][34] = 9'b100000000;
assign Boton[33][35] = 9'b100100000;
assign Boton[33][36] = 9'b100100100;
assign Boton[33][37] = 9'b100000101;
assign Boton[33][38] = 9'b100001001;
assign Boton[33][39] = 9'b100001001;
assign Boton[33][40] = 9'b100101001;
assign Boton[33][41] = 9'b100010011;
assign Boton[33][42] = 9'b100010010;
assign Boton[33][43] = 9'b100000100;
assign Boton[33][44] = 9'b100100100;
assign Boton[34][4] = 9'b100000000;
assign Boton[34][5] = 9'b100100000;
assign Boton[34][6] = 9'b100001001;
assign Boton[34][7] = 9'b100010111;
assign Boton[34][8] = 9'b100001110;
assign Boton[34][9] = 9'b100001001;
assign Boton[34][10] = 9'b100001001;
assign Boton[34][11] = 9'b100000100;
assign Boton[34][12] = 9'b100100100;
assign Boton[34][13] = 9'b100100100;
assign Boton[34][14] = 9'b100000000;
assign Boton[34][15] = 9'b100000000;
assign Boton[34][16] = 9'b100100100;
assign Boton[34][17] = 9'b100000000;
assign Boton[34][18] = 9'b100100000;
assign Boton[34][19] = 9'b100100100;
assign Boton[34][20] = 9'b100001001;
assign Boton[34][21] = 9'b100001001;
assign Boton[34][22] = 9'b100100100;
assign Boton[34][23] = 9'b101101101;
assign Boton[34][24] = 9'b110001101;
assign Boton[34][25] = 9'b110001101;
assign Boton[34][26] = 9'b101101001;
assign Boton[34][27] = 9'b100000100;
assign Boton[34][28] = 9'b100001001;
assign Boton[34][29] = 9'b100100100;
assign Boton[34][30] = 9'b100100100;
assign Boton[34][31] = 9'b100000000;
assign Boton[34][32] = 9'b100000000;
assign Boton[34][33] = 9'b100100100;
assign Boton[34][34] = 9'b100100100;
assign Boton[34][35] = 9'b100100100;
assign Boton[34][36] = 9'b100000000;
assign Boton[34][37] = 9'b100100100;
assign Boton[34][38] = 9'b100001001;
assign Boton[34][39] = 9'b100101001;
assign Boton[34][40] = 9'b100001101;
assign Boton[34][41] = 9'b100011111;
assign Boton[34][42] = 9'b100001101;
assign Boton[34][43] = 9'b100100000;
assign Boton[34][44] = 9'b100000000;
assign Boton[35][4] = 9'b100000000;
assign Boton[35][5] = 9'b100000000;
assign Boton[35][6] = 9'b100100100;
assign Boton[35][7] = 9'b100010010;
assign Boton[35][8] = 9'b100010111;
assign Boton[35][9] = 9'b100001001;
assign Boton[35][10] = 9'b100001001;
assign Boton[35][11] = 9'b100000100;
assign Boton[35][12] = 9'b100000000;
assign Boton[35][13] = 9'b100000000;
assign Boton[35][14] = 9'b100000000;
assign Boton[35][15] = 9'b100000000;
assign Boton[35][16] = 9'b100100100;
assign Boton[35][17] = 9'b100000000;
assign Boton[35][18] = 9'b100000000;
assign Boton[35][19] = 9'b100000000;
assign Boton[35][20] = 9'b100100100;
assign Boton[35][21] = 9'b100101001;
assign Boton[35][22] = 9'b100001001;
assign Boton[35][23] = 9'b100000100;
assign Boton[35][24] = 9'b100000100;
assign Boton[35][25] = 9'b100000100;
assign Boton[35][26] = 9'b100000100;
assign Boton[35][27] = 9'b100000100;
assign Boton[35][28] = 9'b100100100;
assign Boton[35][29] = 9'b100100100;
assign Boton[35][30] = 9'b100100100;
assign Boton[35][31] = 9'b100000000;
assign Boton[35][32] = 9'b100100100;
assign Boton[35][33] = 9'b100100100;
assign Boton[35][34] = 9'b100100100;
assign Boton[35][35] = 9'b100100100;
assign Boton[35][36] = 9'b100100000;
assign Boton[35][37] = 9'b100000100;
assign Boton[35][38] = 9'b100001001;
assign Boton[35][39] = 9'b100001001;
assign Boton[35][40] = 9'b100010010;
assign Boton[35][41] = 9'b100110111;
assign Boton[35][42] = 9'b100100100;
assign Boton[35][43] = 9'b100000000;
assign Boton[35][44] = 9'b100000000;
assign Boton[36][5] = 9'b100000000;
assign Boton[36][6] = 9'b100100000;
assign Boton[36][7] = 9'b100101001;
assign Boton[36][8] = 9'b100010111;
assign Boton[36][9] = 9'b100001101;
assign Boton[36][10] = 9'b100001001;
assign Boton[36][11] = 9'b100000100;
assign Boton[36][12] = 9'b100000000;
assign Boton[36][13] = 9'b100100100;
assign Boton[36][14] = 9'b100100100;
assign Boton[36][15] = 9'b100100100;
assign Boton[36][16] = 9'b100100100;
assign Boton[36][17] = 9'b100000000;
assign Boton[36][18] = 9'b100000000;
assign Boton[36][19] = 9'b100000000;
assign Boton[36][20] = 9'b100000000;
assign Boton[36][21] = 9'b100000000;
assign Boton[36][22] = 9'b100000100;
assign Boton[36][23] = 9'b100001001;
assign Boton[36][24] = 9'b100001001;
assign Boton[36][25] = 9'b100001001;
assign Boton[36][26] = 9'b100000000;
assign Boton[36][27] = 9'b100000000;
assign Boton[36][28] = 9'b100000000;
assign Boton[36][29] = 9'b100000000;
assign Boton[36][30] = 9'b100000000;
assign Boton[36][31] = 9'b100000000;
assign Boton[36][32] = 9'b100000000;
assign Boton[36][33] = 9'b100000000;
assign Boton[36][34] = 9'b100100100;
assign Boton[36][35] = 9'b100100100;
assign Boton[36][36] = 9'b100100000;
assign Boton[36][37] = 9'b100000100;
assign Boton[36][38] = 9'b100001001;
assign Boton[36][39] = 9'b100001101;
assign Boton[36][40] = 9'b100010111;
assign Boton[36][41] = 9'b100101101;
assign Boton[36][42] = 9'b100100000;
assign Boton[36][43] = 9'b100000000;
assign Boton[37][6] = 9'b100000000;
assign Boton[37][7] = 9'b100100100;
assign Boton[37][8] = 9'b100001101;
assign Boton[37][9] = 9'b100010111;
assign Boton[37][10] = 9'b100001001;
assign Boton[37][11] = 9'b100000101;
assign Boton[37][12] = 9'b100000000;
assign Boton[37][13] = 9'b100100100;
assign Boton[37][14] = 9'b100100100;
assign Boton[37][15] = 9'b100100100;
assign Boton[37][16] = 9'b100100100;
assign Boton[37][17] = 9'b101001000;
assign Boton[37][18] = 9'b101101101;
assign Boton[37][19] = 9'b101101101;
assign Boton[37][20] = 9'b101101101;
assign Boton[37][21] = 9'b101101101;
assign Boton[37][22] = 9'b101101101;
assign Boton[37][23] = 9'b101101101;
assign Boton[37][24] = 9'b101110001;
assign Boton[37][25] = 9'b101110001;
assign Boton[37][26] = 9'b101101101;
assign Boton[37][27] = 9'b101101101;
assign Boton[37][28] = 9'b101101101;
assign Boton[37][29] = 9'b101101101;
assign Boton[37][30] = 9'b101101101;
assign Boton[37][31] = 9'b101001000;
assign Boton[37][32] = 9'b100000000;
assign Boton[37][33] = 9'b100000000;
assign Boton[37][34] = 9'b100000000;
assign Boton[37][35] = 9'b100100100;
assign Boton[37][36] = 9'b100100100;
assign Boton[37][37] = 9'b100001001;
assign Boton[37][38] = 9'b100001001;
assign Boton[37][39] = 9'b100010011;
assign Boton[37][40] = 9'b100010010;
assign Boton[37][41] = 9'b100100000;
assign Boton[37][42] = 9'b100100000;
assign Boton[37][43] = 9'b100100100;
assign Boton[38][6] = 9'b100000000;
assign Boton[38][7] = 9'b100100000;
assign Boton[38][8] = 9'b100100100;
assign Boton[38][9] = 9'b100010011;
assign Boton[38][10] = 9'b100010010;
assign Boton[38][11] = 9'b100001001;
assign Boton[38][12] = 9'b100000100;
assign Boton[38][13] = 9'b100100100;
assign Boton[38][14] = 9'b100100100;
assign Boton[38][15] = 9'b100000000;
assign Boton[38][16] = 9'b100100100;
assign Boton[38][17] = 9'b110010001;
assign Boton[38][18] = 9'b111110111;
assign Boton[38][19] = 9'b111110111;
assign Boton[38][20] = 9'b111110111;
assign Boton[38][21] = 9'b111110111;
assign Boton[38][22] = 9'b111110111;
assign Boton[38][23] = 9'b111110111;
assign Boton[38][24] = 9'b111110111;
assign Boton[38][25] = 9'b111110111;
assign Boton[38][26] = 9'b111110111;
assign Boton[38][27] = 9'b111110111;
assign Boton[38][28] = 9'b111110111;
assign Boton[38][29] = 9'b111110111;
assign Boton[38][30] = 9'b111110111;
assign Boton[38][31] = 9'b110110011;
assign Boton[38][32] = 9'b101001000;
assign Boton[38][33] = 9'b100000000;
assign Boton[38][34] = 9'b100100100;
assign Boton[38][35] = 9'b100100100;
assign Boton[38][36] = 9'b100000100;
assign Boton[38][37] = 9'b100001001;
assign Boton[38][38] = 9'b100001110;
assign Boton[38][39] = 9'b100010111;
assign Boton[38][40] = 9'b100100100;
assign Boton[38][41] = 9'b100000000;
assign Boton[38][42] = 9'b100000000;
assign Boton[39][7] = 9'b100000000;
assign Boton[39][8] = 9'b100100000;
assign Boton[39][9] = 9'b100101000;
assign Boton[39][10] = 9'b100010011;
assign Boton[39][11] = 9'b100001101;
assign Boton[39][12] = 9'b100000100;
assign Boton[39][13] = 9'b100100000;
assign Boton[39][14] = 9'b100000000;
assign Boton[39][15] = 9'b100100100;
assign Boton[39][16] = 9'b110010001;
assign Boton[39][17] = 9'b110101111;
assign Boton[39][18] = 9'b101000011;
assign Boton[39][19] = 9'b101000011;
assign Boton[39][20] = 9'b101000011;
assign Boton[39][21] = 9'b101000011;
assign Boton[39][22] = 9'b101000011;
assign Boton[39][23] = 9'b101000011;
assign Boton[39][24] = 9'b101000011;
assign Boton[39][25] = 9'b101000011;
assign Boton[39][26] = 9'b101000011;
assign Boton[39][27] = 9'b101000011;
assign Boton[39][28] = 9'b101000011;
assign Boton[39][29] = 9'b101000011;
assign Boton[39][30] = 9'b101000011;
assign Boton[39][31] = 9'b101100111;
assign Boton[39][32] = 9'b110110011;
assign Boton[39][33] = 9'b100100100;
assign Boton[39][34] = 9'b100100100;
assign Boton[39][35] = 9'b100000100;
assign Boton[39][36] = 9'b100000101;
assign Boton[39][37] = 9'b100001001;
assign Boton[39][38] = 9'b100010011;
assign Boton[39][39] = 9'b100101001;
assign Boton[39][40] = 9'b100100100;
assign Boton[39][41] = 9'b100100100;
assign Boton[40][8] = 9'b100000000;
assign Boton[40][9] = 9'b100100000;
assign Boton[40][10] = 9'b100101000;
assign Boton[40][11] = 9'b100010011;
assign Boton[40][12] = 9'b100001101;
assign Boton[40][13] = 9'b100000000;
assign Boton[40][14] = 9'b100000000;
assign Boton[40][15] = 9'b101101101;
assign Boton[40][16] = 9'b111110111;
assign Boton[40][17] = 9'b101000011;
assign Boton[40][18] = 9'b101000011;
assign Boton[40][19] = 9'b101000011;
assign Boton[40][20] = 9'b101100011;
assign Boton[40][21] = 9'b101100111;
assign Boton[40][22] = 9'b101100011;
assign Boton[40][23] = 9'b101000011;
assign Boton[40][24] = 9'b101000011;
assign Boton[40][25] = 9'b101100011;
assign Boton[40][26] = 9'b101100011;
assign Boton[40][27] = 9'b101100011;
assign Boton[40][28] = 9'b101100011;
assign Boton[40][29] = 9'b101100011;
assign Boton[40][30] = 9'b101000011;
assign Boton[40][31] = 9'b101000011;
assign Boton[40][32] = 9'b110001011;
assign Boton[40][33] = 9'b110110110;
assign Boton[40][34] = 9'b100000000;
assign Boton[40][35] = 9'b100000100;
assign Boton[40][36] = 9'b100001001;
assign Boton[40][37] = 9'b100010011;
assign Boton[40][38] = 9'b100001001;
assign Boton[40][39] = 9'b100100000;
assign Boton[40][40] = 9'b100000000;
assign Boton[41][9] = 9'b100000000;
assign Boton[41][10] = 9'b100000000;
assign Boton[41][11] = 9'b100101000;
assign Boton[41][12] = 9'b100010010;
assign Boton[41][13] = 9'b100001101;
assign Boton[41][14] = 9'b100000000;
assign Boton[41][15] = 9'b101101101;
assign Boton[41][16] = 9'b111110111;
assign Boton[41][17] = 9'b101000011;
assign Boton[41][18] = 9'b101000011;
assign Boton[41][19] = 9'b101100111;
assign Boton[41][20] = 9'b110101111;
assign Boton[41][21] = 9'b101101011;
assign Boton[41][22] = 9'b110001011;
assign Boton[41][23] = 9'b101100111;
assign Boton[41][24] = 9'b110001011;
assign Boton[41][25] = 9'b110001111;
assign Boton[41][26] = 9'b110001111;
assign Boton[41][27] = 9'b110001011;
assign Boton[41][28] = 9'b110110011;
assign Boton[41][29] = 9'b101100111;
assign Boton[41][30] = 9'b101000011;
assign Boton[41][31] = 9'b101000011;
assign Boton[41][32] = 9'b110001011;
assign Boton[41][33] = 9'b110110110;
assign Boton[41][34] = 9'b100000000;
assign Boton[41][35] = 9'b100001001;
assign Boton[41][36] = 9'b100010010;
assign Boton[41][37] = 9'b100101001;
assign Boton[41][38] = 9'b100100000;
assign Boton[41][39] = 9'b100000000;
assign Boton[41][40] = 9'b100000000;
assign Boton[42][10] = 9'b100000000;
assign Boton[42][11] = 9'b100100000;
assign Boton[42][12] = 9'b100101000;
assign Boton[42][13] = 9'b100001101;
assign Boton[42][14] = 9'b100001001;
assign Boton[42][15] = 9'b101001101;
assign Boton[42][16] = 9'b111110011;
assign Boton[42][17] = 9'b101000011;
assign Boton[42][18] = 9'b101000011;
assign Boton[42][19] = 9'b101100111;
assign Boton[42][20] = 9'b110110011;
assign Boton[42][21] = 9'b110001011;
assign Boton[42][22] = 9'b101100011;
assign Boton[42][23] = 9'b110001111;
assign Boton[42][24] = 9'b101100111;
assign Boton[42][25] = 9'b101100111;
assign Boton[42][26] = 9'b101100111;
assign Boton[42][27] = 9'b101000011;
assign Boton[42][28] = 9'b110001011;
assign Boton[42][29] = 9'b101000011;
assign Boton[42][30] = 9'b101000011;
assign Boton[42][31] = 9'b101000011;
assign Boton[42][32] = 9'b110001011;
assign Boton[42][33] = 9'b110010110;
assign Boton[42][34] = 9'b100001001;
assign Boton[42][35] = 9'b100001101;
assign Boton[42][36] = 9'b100000100;
assign Boton[42][37] = 9'b100000000;
assign Boton[42][38] = 9'b100000000;
assign Boton[42][39] = 9'b100000100;
assign Boton[43][11] = 9'b100000000;
assign Boton[43][12] = 9'b100100000;
assign Boton[43][13] = 9'b100100100;
assign Boton[43][14] = 9'b100001001;
assign Boton[43][15] = 9'b101110001;
assign Boton[43][16] = 9'b111110011;
assign Boton[43][17] = 9'b101000011;
assign Boton[43][18] = 9'b101000011;
assign Boton[43][19] = 9'b101100111;
assign Boton[43][20] = 9'b110110011;
assign Boton[43][21] = 9'b101101011;
assign Boton[43][22] = 9'b110001011;
assign Boton[43][23] = 9'b110001011;
assign Boton[43][24] = 9'b110001011;
assign Boton[43][25] = 9'b110001111;
assign Boton[43][26] = 9'b110001011;
assign Boton[43][27] = 9'b101100011;
assign Boton[43][28] = 9'b110001111;
assign Boton[43][29] = 9'b101000011;
assign Boton[43][30] = 9'b101000011;
assign Boton[43][31] = 9'b101000011;
assign Boton[43][32] = 9'b110001011;
assign Boton[43][33] = 9'b110011111;
assign Boton[43][34] = 9'b100001001;
assign Boton[43][35] = 9'b100100100;
assign Boton[43][36] = 9'b100100000;
assign Boton[43][37] = 9'b100000000;
assign Boton[44][12] = 9'b100000000;
assign Boton[44][13] = 9'b100000000;
assign Boton[44][14] = 9'b100000000;
assign Boton[44][15] = 9'b101101101;
assign Boton[44][16] = 9'b111110111;
assign Boton[44][17] = 9'b101000011;
assign Boton[44][18] = 9'b101000011;
assign Boton[44][19] = 9'b101100011;
assign Boton[44][20] = 9'b110001011;
assign Boton[44][21] = 9'b110001011;
assign Boton[44][22] = 9'b101100111;
assign Boton[44][23] = 9'b101000011;
assign Boton[44][24] = 9'b101100011;
assign Boton[44][25] = 9'b110001011;
assign Boton[44][26] = 9'b110001011;
assign Boton[44][27] = 9'b101000011;
assign Boton[44][28] = 9'b101100111;
assign Boton[44][29] = 9'b101000011;
assign Boton[44][30] = 9'b101000011;
assign Boton[44][31] = 9'b101000011;
assign Boton[44][32] = 9'b110001011;
assign Boton[44][33] = 9'b110111110;
assign Boton[44][34] = 9'b100000000;
assign Boton[44][35] = 9'b100100100;
assign Boton[44][36] = 9'b100100100;
assign Boton[45][13] = 9'b100000000;
assign Boton[45][14] = 9'b100000000;
assign Boton[45][15] = 9'b100101000;
assign Boton[45][16] = 9'b110010010;
assign Boton[45][17] = 9'b110001011;
assign Boton[45][18] = 9'b101000011;
assign Boton[45][19] = 9'b101000011;
assign Boton[45][20] = 9'b101000011;
assign Boton[45][21] = 9'b101000011;
assign Boton[45][22] = 9'b101000011;
assign Boton[45][23] = 9'b101000011;
assign Boton[45][24] = 9'b101000011;
assign Boton[45][25] = 9'b101000011;
assign Boton[45][26] = 9'b101000011;
assign Boton[45][27] = 9'b101100011;
assign Boton[45][28] = 9'b101000011;
assign Boton[45][29] = 9'b101100011;
assign Boton[45][30] = 9'b101000011;
assign Boton[45][31] = 9'b101100111;
assign Boton[45][32] = 9'b110110011;
assign Boton[45][33] = 9'b101101101;
assign Boton[45][34] = 9'b100000000;
assign Boton[45][35] = 9'b100100100;
assign Boton[46][15] = 9'b100000000;
assign Boton[46][16] = 9'b101001000;
assign Boton[46][17] = 9'b110010010;
assign Boton[46][18] = 9'b101000011;
assign Boton[46][19] = 9'b101000011;
assign Boton[46][20] = 9'b101000011;
assign Boton[46][21] = 9'b101000011;
assign Boton[46][22] = 9'b101100011;
assign Boton[46][23] = 9'b101100011;
assign Boton[46][24] = 9'b110001011;
assign Boton[46][25] = 9'b101100111;
assign Boton[46][26] = 9'b101100011;
assign Boton[46][27] = 9'b101000011;
assign Boton[46][28] = 9'b101000011;
assign Boton[46][29] = 9'b101000011;
assign Boton[46][30] = 9'b101000011;
assign Boton[46][31] = 9'b110001011;
assign Boton[46][32] = 9'b101110001;
assign Boton[46][33] = 9'b100000000;
assign Boton[47][22] = 9'b101101101;
assign Boton[47][23] = 9'b110110110;
assign Boton[47][24] = 9'b111111111;
assign Boton[47][25] = 9'b111111111;
assign Boton[47][26] = 9'b111111110;
//Total de Lineas = 1667
endmodule

